`timescale 1ns / 1ps

module lut_exp_19in_16out(
    input  signed [18:0] in,
    output        [15:0] exp
    );
    
    reg  [18:0] addr;
    reg  [15:0] exp_inner;
    reg  [15:0] exp_table[0:2047];
    initial begin
exp_table[11'b10000000000] = 16'b0000000100101100;
	exp_table[11'b10000000001] = 16'b0000000100101101;
	exp_table[11'b10000000010] = 16'b0000000100101110;
	exp_table[11'b10000000011] = 16'b0000000100101111;
	exp_table[11'b10000000100] = 16'b0000000100110000;
	exp_table[11'b10000000101] = 16'b0000000100110010;
	exp_table[11'b10000000110] = 16'b0000000100110011;
	exp_table[11'b10000000111] = 16'b0000000100110100;
	exp_table[11'b10000001000] = 16'b0000000100110101;
	exp_table[11'b10000001001] = 16'b0000000100110110;
	exp_table[11'b10000001010] = 16'b0000000100111000;
	exp_table[11'b10000001011] = 16'b0000000100111001;
	exp_table[11'b10000001100] = 16'b0000000100111010;
	exp_table[11'b10000001101] = 16'b0000000100111011;
	exp_table[11'b10000001110] = 16'b0000000100111100;
	exp_table[11'b10000001111] = 16'b0000000100111110;
	exp_table[11'b10000010000] = 16'b0000000100111111;
	exp_table[11'b10000010001] = 16'b0000000101000000;
	exp_table[11'b10000010010] = 16'b0000000101000001;
	exp_table[11'b10000010011] = 16'b0000000101000011;
	exp_table[11'b10000010100] = 16'b0000000101000100;
	exp_table[11'b10000010101] = 16'b0000000101000101;
	exp_table[11'b10000010110] = 16'b0000000101000111;
	exp_table[11'b10000010111] = 16'b0000000101001000;
	exp_table[11'b10000011000] = 16'b0000000101001001;
	exp_table[11'b10000011001] = 16'b0000000101001010;
	exp_table[11'b10000011010] = 16'b0000000101001100;
	exp_table[11'b10000011011] = 16'b0000000101001101;
	exp_table[11'b10000011100] = 16'b0000000101001110;
	exp_table[11'b10000011101] = 16'b0000000101010000;
	exp_table[11'b10000011110] = 16'b0000000101010001;
	exp_table[11'b10000011111] = 16'b0000000101010010;
	exp_table[11'b10000100000] = 16'b0000000101010100;
	exp_table[11'b10000100001] = 16'b0000000101010101;
	exp_table[11'b10000100010] = 16'b0000000101010110;
	exp_table[11'b10000100011] = 16'b0000000101011000;
	exp_table[11'b10000100100] = 16'b0000000101011001;
	exp_table[11'b10000100101] = 16'b0000000101011010;
	exp_table[11'b10000100110] = 16'b0000000101011100;
	exp_table[11'b10000100111] = 16'b0000000101011101;
	exp_table[11'b10000101000] = 16'b0000000101011110;
	exp_table[11'b10000101001] = 16'b0000000101100000;
	exp_table[11'b10000101010] = 16'b0000000101100001;
	exp_table[11'b10000101011] = 16'b0000000101100010;
	exp_table[11'b10000101100] = 16'b0000000101100100;
	exp_table[11'b10000101101] = 16'b0000000101100101;
	exp_table[11'b10000101110] = 16'b0000000101100111;
	exp_table[11'b10000101111] = 16'b0000000101101000;
	exp_table[11'b10000110000] = 16'b0000000101101001;
	exp_table[11'b10000110001] = 16'b0000000101101011;
	exp_table[11'b10000110010] = 16'b0000000101101100;
	exp_table[11'b10000110011] = 16'b0000000101101110;
	exp_table[11'b10000110100] = 16'b0000000101101111;
	exp_table[11'b10000110101] = 16'b0000000101110001;
	exp_table[11'b10000110110] = 16'b0000000101110010;
	exp_table[11'b10000110111] = 16'b0000000101110100;
	exp_table[11'b10000111000] = 16'b0000000101110101;
	exp_table[11'b10000111001] = 16'b0000000101110110;
	exp_table[11'b10000111010] = 16'b0000000101111000;
	exp_table[11'b10000111011] = 16'b0000000101111001;
	exp_table[11'b10000111100] = 16'b0000000101111011;
	exp_table[11'b10000111101] = 16'b0000000101111100;
	exp_table[11'b10000111110] = 16'b0000000101111110;
	exp_table[11'b10000111111] = 16'b0000000101111111;
	exp_table[11'b10001000000] = 16'b0000000110000001;
	exp_table[11'b10001000001] = 16'b0000000110000010;
	exp_table[11'b10001000010] = 16'b0000000110000100;
	exp_table[11'b10001000011] = 16'b0000000110000101;
	exp_table[11'b10001000100] = 16'b0000000110000111;
	exp_table[11'b10001000101] = 16'b0000000110001000;
	exp_table[11'b10001000110] = 16'b0000000110001010;
	exp_table[11'b10001000111] = 16'b0000000110001011;
	exp_table[11'b10001001000] = 16'b0000000110001101;
	exp_table[11'b10001001001] = 16'b0000000110001111;
	exp_table[11'b10001001010] = 16'b0000000110010000;
	exp_table[11'b10001001011] = 16'b0000000110010010;
	exp_table[11'b10001001100] = 16'b0000000110010011;
	exp_table[11'b10001001101] = 16'b0000000110010101;
	exp_table[11'b10001001110] = 16'b0000000110010110;
	exp_table[11'b10001001111] = 16'b0000000110011000;
	exp_table[11'b10001010000] = 16'b0000000110011010;
	exp_table[11'b10001010001] = 16'b0000000110011011;
	exp_table[11'b10001010010] = 16'b0000000110011101;
	exp_table[11'b10001010011] = 16'b0000000110011111;
	exp_table[11'b10001010100] = 16'b0000000110100000;
	exp_table[11'b10001010101] = 16'b0000000110100010;
	exp_table[11'b10001010110] = 16'b0000000110100011;
	exp_table[11'b10001010111] = 16'b0000000110100101;
	exp_table[11'b10001011000] = 16'b0000000110100111;
	exp_table[11'b10001011001] = 16'b0000000110101000;
	exp_table[11'b10001011010] = 16'b0000000110101010;
	exp_table[11'b10001011011] = 16'b0000000110101100;
	exp_table[11'b10001011100] = 16'b0000000110101101;
	exp_table[11'b10001011101] = 16'b0000000110101111;
	exp_table[11'b10001011110] = 16'b0000000110110001;
	exp_table[11'b10001011111] = 16'b0000000110110010;
	exp_table[11'b10001100000] = 16'b0000000110110100;
	exp_table[11'b10001100001] = 16'b0000000110110110;
	exp_table[11'b10001100010] = 16'b0000000110111000;
	exp_table[11'b10001100011] = 16'b0000000110111001;
	exp_table[11'b10001100100] = 16'b0000000110111011;
	exp_table[11'b10001100101] = 16'b0000000110111101;
	exp_table[11'b10001100110] = 16'b0000000110111110;
	exp_table[11'b10001100111] = 16'b0000000111000000;
	exp_table[11'b10001101000] = 16'b0000000111000010;
	exp_table[11'b10001101001] = 16'b0000000111000100;
	exp_table[11'b10001101010] = 16'b0000000111000110;
	exp_table[11'b10001101011] = 16'b0000000111000111;
	exp_table[11'b10001101100] = 16'b0000000111001001;
	exp_table[11'b10001101101] = 16'b0000000111001011;
	exp_table[11'b10001101110] = 16'b0000000111001101;
	exp_table[11'b10001101111] = 16'b0000000111001110;
	exp_table[11'b10001110000] = 16'b0000000111010000;
	exp_table[11'b10001110001] = 16'b0000000111010010;
	exp_table[11'b10001110010] = 16'b0000000111010100;
	exp_table[11'b10001110011] = 16'b0000000111010110;
	exp_table[11'b10001110100] = 16'b0000000111011000;
	exp_table[11'b10001110101] = 16'b0000000111011001;
	exp_table[11'b10001110110] = 16'b0000000111011011;
	exp_table[11'b10001110111] = 16'b0000000111011101;
	exp_table[11'b10001111000] = 16'b0000000111011111;
	exp_table[11'b10001111001] = 16'b0000000111100001;
	exp_table[11'b10001111010] = 16'b0000000111100011;
	exp_table[11'b10001111011] = 16'b0000000111100101;
	exp_table[11'b10001111100] = 16'b0000000111100111;
	exp_table[11'b10001111101] = 16'b0000000111101000;
	exp_table[11'b10001111110] = 16'b0000000111101010;
	exp_table[11'b10001111111] = 16'b0000000111101100;
	exp_table[11'b10010000000] = 16'b0000000111101110;
	exp_table[11'b10010000001] = 16'b0000000111110000;
	exp_table[11'b10010000010] = 16'b0000000111110010;
	exp_table[11'b10010000011] = 16'b0000000111110100;
	exp_table[11'b10010000100] = 16'b0000000111110110;
	exp_table[11'b10010000101] = 16'b0000000111111000;
	exp_table[11'b10010000110] = 16'b0000000111111010;
	exp_table[11'b10010000111] = 16'b0000000111111100;
	exp_table[11'b10010001000] = 16'b0000000111111110;
	exp_table[11'b10010001001] = 16'b0000001000000000;
	exp_table[11'b10010001010] = 16'b0000001000000010;
	exp_table[11'b10010001011] = 16'b0000001000000100;
	exp_table[11'b10010001100] = 16'b0000001000000110;
	exp_table[11'b10010001101] = 16'b0000001000001000;
	exp_table[11'b10010001110] = 16'b0000001000001010;
	exp_table[11'b10010001111] = 16'b0000001000001100;
	exp_table[11'b10010010000] = 16'b0000001000001110;
	exp_table[11'b10010010001] = 16'b0000001000010000;
	exp_table[11'b10010010010] = 16'b0000001000010010;
	exp_table[11'b10010010011] = 16'b0000001000010100;
	exp_table[11'b10010010100] = 16'b0000001000010110;
	exp_table[11'b10010010101] = 16'b0000001000011001;
	exp_table[11'b10010010110] = 16'b0000001000011011;
	exp_table[11'b10010010111] = 16'b0000001000011101;
	exp_table[11'b10010011000] = 16'b0000001000011111;
	exp_table[11'b10010011001] = 16'b0000001000100001;
	exp_table[11'b10010011010] = 16'b0000001000100011;
	exp_table[11'b10010011011] = 16'b0000001000100101;
	exp_table[11'b10010011100] = 16'b0000001000100111;
	exp_table[11'b10010011101] = 16'b0000001000101010;
	exp_table[11'b10010011110] = 16'b0000001000101100;
	exp_table[11'b10010011111] = 16'b0000001000101110;
	exp_table[11'b10010100000] = 16'b0000001000110000;
	exp_table[11'b10010100001] = 16'b0000001000110010;
	exp_table[11'b10010100010] = 16'b0000001000110101;
	exp_table[11'b10010100011] = 16'b0000001000110111;
	exp_table[11'b10010100100] = 16'b0000001000111001;
	exp_table[11'b10010100101] = 16'b0000001000111011;
	exp_table[11'b10010100110] = 16'b0000001000111101;
	exp_table[11'b10010100111] = 16'b0000001001000000;
	exp_table[11'b10010101000] = 16'b0000001001000010;
	exp_table[11'b10010101001] = 16'b0000001001000100;
	exp_table[11'b10010101010] = 16'b0000001001000110;
	exp_table[11'b10010101011] = 16'b0000001001001001;
	exp_table[11'b10010101100] = 16'b0000001001001011;
	exp_table[11'b10010101101] = 16'b0000001001001101;
	exp_table[11'b10010101110] = 16'b0000001001010000;
	exp_table[11'b10010101111] = 16'b0000001001010010;
	exp_table[11'b10010110000] = 16'b0000001001010100;
	exp_table[11'b10010110001] = 16'b0000001001010111;
	exp_table[11'b10010110010] = 16'b0000001001011001;
	exp_table[11'b10010110011] = 16'b0000001001011011;
	exp_table[11'b10010110100] = 16'b0000001001011110;
	exp_table[11'b10010110101] = 16'b0000001001100000;
	exp_table[11'b10010110110] = 16'b0000001001100010;
	exp_table[11'b10010110111] = 16'b0000001001100101;
	exp_table[11'b10010111000] = 16'b0000001001100111;
	exp_table[11'b10010111001] = 16'b0000001001101010;
	exp_table[11'b10010111010] = 16'b0000001001101100;
	exp_table[11'b10010111011] = 16'b0000001001101110;
	exp_table[11'b10010111100] = 16'b0000001001110001;
	exp_table[11'b10010111101] = 16'b0000001001110011;
	exp_table[11'b10010111110] = 16'b0000001001110110;
	exp_table[11'b10010111111] = 16'b0000001001111000;
	exp_table[11'b10011000000] = 16'b0000001001111011;
	exp_table[11'b10011000001] = 16'b0000001001111101;
	exp_table[11'b10011000010] = 16'b0000001010000000;
	exp_table[11'b10011000011] = 16'b0000001010000010;
	exp_table[11'b10011000100] = 16'b0000001010000101;
	exp_table[11'b10011000101] = 16'b0000001010000111;
	exp_table[11'b10011000110] = 16'b0000001010001010;
	exp_table[11'b10011000111] = 16'b0000001010001100;
	exp_table[11'b10011001000] = 16'b0000001010001111;
	exp_table[11'b10011001001] = 16'b0000001010010010;
	exp_table[11'b10011001010] = 16'b0000001010010100;
	exp_table[11'b10011001011] = 16'b0000001010010111;
	exp_table[11'b10011001100] = 16'b0000001010011001;
	exp_table[11'b10011001101] = 16'b0000001010011100;
	exp_table[11'b10011001110] = 16'b0000001010011110;
	exp_table[11'b10011001111] = 16'b0000001010100001;
	exp_table[11'b10011010000] = 16'b0000001010100100;
	exp_table[11'b10011010001] = 16'b0000001010100110;
	exp_table[11'b10011010010] = 16'b0000001010101001;
	exp_table[11'b10011010011] = 16'b0000001010101100;
	exp_table[11'b10011010100] = 16'b0000001010101110;
	exp_table[11'b10011010101] = 16'b0000001010110001;
	exp_table[11'b10011010110] = 16'b0000001010110100;
	exp_table[11'b10011010111] = 16'b0000001010110110;
	exp_table[11'b10011011000] = 16'b0000001010111001;
	exp_table[11'b10011011001] = 16'b0000001010111100;
	exp_table[11'b10011011010] = 16'b0000001010111111;
	exp_table[11'b10011011011] = 16'b0000001011000001;
	exp_table[11'b10011011100] = 16'b0000001011000100;
	exp_table[11'b10011011101] = 16'b0000001011000111;
	exp_table[11'b10011011110] = 16'b0000001011001010;
	exp_table[11'b10011011111] = 16'b0000001011001101;
	exp_table[11'b10011100000] = 16'b0000001011001111;
	exp_table[11'b10011100001] = 16'b0000001011010010;
	exp_table[11'b10011100010] = 16'b0000001011010101;
	exp_table[11'b10011100011] = 16'b0000001011011000;
	exp_table[11'b10011100100] = 16'b0000001011011011;
	exp_table[11'b10011100101] = 16'b0000001011011110;
	exp_table[11'b10011100110] = 16'b0000001011100000;
	exp_table[11'b10011100111] = 16'b0000001011100011;
	exp_table[11'b10011101000] = 16'b0000001011100110;
	exp_table[11'b10011101001] = 16'b0000001011101001;
	exp_table[11'b10011101010] = 16'b0000001011101100;
	exp_table[11'b10011101011] = 16'b0000001011101111;
	exp_table[11'b10011101100] = 16'b0000001011110010;
	exp_table[11'b10011101101] = 16'b0000001011110101;
	exp_table[11'b10011101110] = 16'b0000001011111000;
	exp_table[11'b10011101111] = 16'b0000001011111011;
	exp_table[11'b10011110000] = 16'b0000001011111110;
	exp_table[11'b10011110001] = 16'b0000001100000001;
	exp_table[11'b10011110010] = 16'b0000001100000100;
	exp_table[11'b10011110011] = 16'b0000001100000111;
	exp_table[11'b10011110100] = 16'b0000001100001010;
	exp_table[11'b10011110101] = 16'b0000001100001101;
	exp_table[11'b10011110110] = 16'b0000001100010000;
	exp_table[11'b10011110111] = 16'b0000001100010011;
	exp_table[11'b10011111000] = 16'b0000001100010110;
	exp_table[11'b10011111001] = 16'b0000001100011001;
	exp_table[11'b10011111010] = 16'b0000001100011100;
	exp_table[11'b10011111011] = 16'b0000001100011111;
	exp_table[11'b10011111100] = 16'b0000001100100011;
	exp_table[11'b10011111101] = 16'b0000001100100110;
	exp_table[11'b10011111110] = 16'b0000001100101001;
	exp_table[11'b10011111111] = 16'b0000001100101100;
	exp_table[11'b10100000000] = 16'b0000001100101111;
	exp_table[11'b10100000001] = 16'b0000001100110010;
	exp_table[11'b10100000010] = 16'b0000001100110110;
	exp_table[11'b10100000011] = 16'b0000001100111001;
	exp_table[11'b10100000100] = 16'b0000001100111100;
	exp_table[11'b10100000101] = 16'b0000001100111111;
	exp_table[11'b10100000110] = 16'b0000001101000011;
	exp_table[11'b10100000111] = 16'b0000001101000110;
	exp_table[11'b10100001000] = 16'b0000001101001001;
	exp_table[11'b10100001001] = 16'b0000001101001100;
	exp_table[11'b10100001010] = 16'b0000001101010000;
	exp_table[11'b10100001011] = 16'b0000001101010011;
	exp_table[11'b10100001100] = 16'b0000001101010110;
	exp_table[11'b10100001101] = 16'b0000001101011010;
	exp_table[11'b10100001110] = 16'b0000001101011101;
	exp_table[11'b10100001111] = 16'b0000001101100000;
	exp_table[11'b10100010000] = 16'b0000001101100100;
	exp_table[11'b10100010001] = 16'b0000001101100111;
	exp_table[11'b10100010010] = 16'b0000001101101011;
	exp_table[11'b10100010011] = 16'b0000001101101110;
	exp_table[11'b10100010100] = 16'b0000001101110001;
	exp_table[11'b10100010101] = 16'b0000001101110101;
	exp_table[11'b10100010110] = 16'b0000001101111000;
	exp_table[11'b10100010111] = 16'b0000001101111100;
	exp_table[11'b10100011000] = 16'b0000001101111111;
	exp_table[11'b10100011001] = 16'b0000001110000011;
	exp_table[11'b10100011010] = 16'b0000001110000110;
	exp_table[11'b10100011011] = 16'b0000001110001010;
	exp_table[11'b10100011100] = 16'b0000001110001101;
	exp_table[11'b10100011101] = 16'b0000001110010001;
	exp_table[11'b10100011110] = 16'b0000001110010101;
	exp_table[11'b10100011111] = 16'b0000001110011000;
	exp_table[11'b10100100000] = 16'b0000001110011100;
	exp_table[11'b10100100001] = 16'b0000001110011111;
	exp_table[11'b10100100010] = 16'b0000001110100011;
	exp_table[11'b10100100011] = 16'b0000001110100111;
	exp_table[11'b10100100100] = 16'b0000001110101010;
	exp_table[11'b10100100101] = 16'b0000001110101110;
	exp_table[11'b10100100110] = 16'b0000001110110010;
	exp_table[11'b10100100111] = 16'b0000001110110101;
	exp_table[11'b10100101000] = 16'b0000001110111001;
	exp_table[11'b10100101001] = 16'b0000001110111101;
	exp_table[11'b10100101010] = 16'b0000001111000001;
	exp_table[11'b10100101011] = 16'b0000001111000100;
	exp_table[11'b10100101100] = 16'b0000001111001000;
	exp_table[11'b10100101101] = 16'b0000001111001100;
	exp_table[11'b10100101110] = 16'b0000001111010000;
	exp_table[11'b10100101111] = 16'b0000001111010100;
	exp_table[11'b10100110000] = 16'b0000001111010111;
	exp_table[11'b10100110001] = 16'b0000001111011011;
	exp_table[11'b10100110010] = 16'b0000001111011111;
	exp_table[11'b10100110011] = 16'b0000001111100011;
	exp_table[11'b10100110100] = 16'b0000001111100111;
	exp_table[11'b10100110101] = 16'b0000001111101011;
	exp_table[11'b10100110110] = 16'b0000001111101111;
	exp_table[11'b10100110111] = 16'b0000001111110011;
	exp_table[11'b10100111000] = 16'b0000001111110111;
	exp_table[11'b10100111001] = 16'b0000001111111011;
	exp_table[11'b10100111010] = 16'b0000001111111111;
	exp_table[11'b10100111011] = 16'b0000010000000011;
	exp_table[11'b10100111100] = 16'b0000010000000111;
	exp_table[11'b10100111101] = 16'b0000010000001011;
	exp_table[11'b10100111110] = 16'b0000010000001111;
	exp_table[11'b10100111111] = 16'b0000010000010011;
	exp_table[11'b10101000000] = 16'b0000010000010111;
	exp_table[11'b10101000001] = 16'b0000010000011011;
	exp_table[11'b10101000010] = 16'b0000010000011111;
	exp_table[11'b10101000011] = 16'b0000010000100011;
	exp_table[11'b10101000100] = 16'b0000010000100111;
	exp_table[11'b10101000101] = 16'b0000010000101100;
	exp_table[11'b10101000110] = 16'b0000010000110000;
	exp_table[11'b10101000111] = 16'b0000010000110100;
	exp_table[11'b10101001000] = 16'b0000010000111000;
	exp_table[11'b10101001001] = 16'b0000010000111100;
	exp_table[11'b10101001010] = 16'b0000010001000001;
	exp_table[11'b10101001011] = 16'b0000010001000101;
	exp_table[11'b10101001100] = 16'b0000010001001001;
	exp_table[11'b10101001101] = 16'b0000010001001101;
	exp_table[11'b10101001110] = 16'b0000010001010010;
	exp_table[11'b10101001111] = 16'b0000010001010110;
	exp_table[11'b10101010000] = 16'b0000010001011010;
	exp_table[11'b10101010001] = 16'b0000010001011111;
	exp_table[11'b10101010010] = 16'b0000010001100011;
	exp_table[11'b10101010011] = 16'b0000010001101000;
	exp_table[11'b10101010100] = 16'b0000010001101100;
	exp_table[11'b10101010101] = 16'b0000010001110000;
	exp_table[11'b10101010110] = 16'b0000010001110101;
	exp_table[11'b10101010111] = 16'b0000010001111001;
	exp_table[11'b10101011000] = 16'b0000010001111110;
	exp_table[11'b10101011001] = 16'b0000010010000010;
	exp_table[11'b10101011010] = 16'b0000010010000111;
	exp_table[11'b10101011011] = 16'b0000010010001011;
	exp_table[11'b10101011100] = 16'b0000010010010000;
	exp_table[11'b10101011101] = 16'b0000010010010101;
	exp_table[11'b10101011110] = 16'b0000010010011001;
	exp_table[11'b10101011111] = 16'b0000010010011110;
	exp_table[11'b10101100000] = 16'b0000010010100010;
	exp_table[11'b10101100001] = 16'b0000010010100111;
	exp_table[11'b10101100010] = 16'b0000010010101100;
	exp_table[11'b10101100011] = 16'b0000010010110000;
	exp_table[11'b10101100100] = 16'b0000010010110101;
	exp_table[11'b10101100101] = 16'b0000010010111010;
	exp_table[11'b10101100110] = 16'b0000010010111110;
	exp_table[11'b10101100111] = 16'b0000010011000011;
	exp_table[11'b10101101000] = 16'b0000010011001000;
	exp_table[11'b10101101001] = 16'b0000010011001101;
	exp_table[11'b10101101010] = 16'b0000010011010010;
	exp_table[11'b10101101011] = 16'b0000010011010110;
	exp_table[11'b10101101100] = 16'b0000010011011011;
	exp_table[11'b10101101101] = 16'b0000010011100000;
	exp_table[11'b10101101110] = 16'b0000010011100101;
	exp_table[11'b10101101111] = 16'b0000010011101010;
	exp_table[11'b10101110000] = 16'b0000010011101111;
	exp_table[11'b10101110001] = 16'b0000010011110100;
	exp_table[11'b10101110010] = 16'b0000010011111001;
	exp_table[11'b10101110011] = 16'b0000010011111110;
	exp_table[11'b10101110100] = 16'b0000010100000011;
	exp_table[11'b10101110101] = 16'b0000010100001000;
	exp_table[11'b10101110110] = 16'b0000010100001101;
	exp_table[11'b10101110111] = 16'b0000010100010010;
	exp_table[11'b10101111000] = 16'b0000010100010111;
	exp_table[11'b10101111001] = 16'b0000010100011100;
	exp_table[11'b10101111010] = 16'b0000010100100001;
	exp_table[11'b10101111011] = 16'b0000010100100110;
	exp_table[11'b10101111100] = 16'b0000010100101100;
	exp_table[11'b10101111101] = 16'b0000010100110001;
	exp_table[11'b10101111110] = 16'b0000010100110110;
	exp_table[11'b10101111111] = 16'b0000010100111011;
	exp_table[11'b10110000000] = 16'b0000010101000000;
	exp_table[11'b10110000001] = 16'b0000010101000110;
	exp_table[11'b10110000010] = 16'b0000010101001011;
	exp_table[11'b10110000011] = 16'b0000010101010000;
	exp_table[11'b10110000100] = 16'b0000010101010110;
	exp_table[11'b10110000101] = 16'b0000010101011011;
	exp_table[11'b10110000110] = 16'b0000010101100000;
	exp_table[11'b10110000111] = 16'b0000010101100110;
	exp_table[11'b10110001000] = 16'b0000010101101011;
	exp_table[11'b10110001001] = 16'b0000010101110001;
	exp_table[11'b10110001010] = 16'b0000010101110110;
	exp_table[11'b10110001011] = 16'b0000010101111011;
	exp_table[11'b10110001100] = 16'b0000010110000001;
	exp_table[11'b10110001101] = 16'b0000010110000110;
	exp_table[11'b10110001110] = 16'b0000010110001100;
	exp_table[11'b10110001111] = 16'b0000010110010010;
	exp_table[11'b10110010000] = 16'b0000010110010111;
	exp_table[11'b10110010001] = 16'b0000010110011101;
	exp_table[11'b10110010010] = 16'b0000010110100010;
	exp_table[11'b10110010011] = 16'b0000010110101000;
	exp_table[11'b10110010100] = 16'b0000010110101110;
	exp_table[11'b10110010101] = 16'b0000010110110011;
	exp_table[11'b10110010110] = 16'b0000010110111001;
	exp_table[11'b10110010111] = 16'b0000010110111111;
	exp_table[11'b10110011000] = 16'b0000010111000101;
	exp_table[11'b10110011001] = 16'b0000010111001010;
	exp_table[11'b10110011010] = 16'b0000010111010000;
	exp_table[11'b10110011011] = 16'b0000010111010110;
	exp_table[11'b10110011100] = 16'b0000010111011100;
	exp_table[11'b10110011101] = 16'b0000010111100010;
	exp_table[11'b10110011110] = 16'b0000010111101000;
	exp_table[11'b10110011111] = 16'b0000010111101110;
	exp_table[11'b10110100000] = 16'b0000010111110011;
	exp_table[11'b10110100001] = 16'b0000010111111001;
	exp_table[11'b10110100010] = 16'b0000010111111111;
	exp_table[11'b10110100011] = 16'b0000011000000101;
	exp_table[11'b10110100100] = 16'b0000011000001011;
	exp_table[11'b10110100101] = 16'b0000011000010010;
	exp_table[11'b10110100110] = 16'b0000011000011000;
	exp_table[11'b10110100111] = 16'b0000011000011110;
	exp_table[11'b10110101000] = 16'b0000011000100100;
	exp_table[11'b10110101001] = 16'b0000011000101010;
	exp_table[11'b10110101010] = 16'b0000011000110000;
	exp_table[11'b10110101011] = 16'b0000011000110110;
	exp_table[11'b10110101100] = 16'b0000011000111101;
	exp_table[11'b10110101101] = 16'b0000011001000011;
	exp_table[11'b10110101110] = 16'b0000011001001001;
	exp_table[11'b10110101111] = 16'b0000011001001111;
	exp_table[11'b10110110000] = 16'b0000011001010110;
	exp_table[11'b10110110001] = 16'b0000011001011100;
	exp_table[11'b10110110010] = 16'b0000011001100010;
	exp_table[11'b10110110011] = 16'b0000011001101001;
	exp_table[11'b10110110100] = 16'b0000011001101111;
	exp_table[11'b10110110101] = 16'b0000011001110110;
	exp_table[11'b10110110110] = 16'b0000011001111100;
	exp_table[11'b10110110111] = 16'b0000011010000011;
	exp_table[11'b10110111000] = 16'b0000011010001001;
	exp_table[11'b10110111001] = 16'b0000011010010000;
	exp_table[11'b10110111010] = 16'b0000011010010110;
	exp_table[11'b10110111011] = 16'b0000011010011101;
	exp_table[11'b10110111100] = 16'b0000011010100100;
	exp_table[11'b10110111101] = 16'b0000011010101010;
	exp_table[11'b10110111110] = 16'b0000011010110001;
	exp_table[11'b10110111111] = 16'b0000011010111000;
	exp_table[11'b10111000000] = 16'b0000011010111110;
	exp_table[11'b10111000001] = 16'b0000011011000101;
	exp_table[11'b10111000010] = 16'b0000011011001100;
	exp_table[11'b10111000011] = 16'b0000011011010011;
	exp_table[11'b10111000100] = 16'b0000011011011010;
	exp_table[11'b10111000101] = 16'b0000011011100000;
	exp_table[11'b10111000110] = 16'b0000011011100111;
	exp_table[11'b10111000111] = 16'b0000011011101110;
	exp_table[11'b10111001000] = 16'b0000011011110101;
	exp_table[11'b10111001001] = 16'b0000011011111100;
	exp_table[11'b10111001010] = 16'b0000011100000011;
	exp_table[11'b10111001011] = 16'b0000011100001010;
	exp_table[11'b10111001100] = 16'b0000011100010001;
	exp_table[11'b10111001101] = 16'b0000011100011000;
	exp_table[11'b10111001110] = 16'b0000011100011111;
	exp_table[11'b10111001111] = 16'b0000011100100111;
	exp_table[11'b10111010000] = 16'b0000011100101110;
	exp_table[11'b10111010001] = 16'b0000011100110101;
	exp_table[11'b10111010010] = 16'b0000011100111100;
	exp_table[11'b10111010011] = 16'b0000011101000011;
	exp_table[11'b10111010100] = 16'b0000011101001011;
	exp_table[11'b10111010101] = 16'b0000011101010010;
	exp_table[11'b10111010110] = 16'b0000011101011001;
	exp_table[11'b10111010111] = 16'b0000011101100001;
	exp_table[11'b10111011000] = 16'b0000011101101000;
	exp_table[11'b10111011001] = 16'b0000011101110000;
	exp_table[11'b10111011010] = 16'b0000011101110111;
	exp_table[11'b10111011011] = 16'b0000011101111110;
	exp_table[11'b10111011100] = 16'b0000011110000110;
	exp_table[11'b10111011101] = 16'b0000011110001101;
	exp_table[11'b10111011110] = 16'b0000011110010101;
	exp_table[11'b10111011111] = 16'b0000011110011101;
	exp_table[11'b10111100000] = 16'b0000011110100100;
	exp_table[11'b10111100001] = 16'b0000011110101100;
	exp_table[11'b10111100010] = 16'b0000011110110100;
	exp_table[11'b10111100011] = 16'b0000011110111011;
	exp_table[11'b10111100100] = 16'b0000011111000011;
	exp_table[11'b10111100101] = 16'b0000011111001011;
	exp_table[11'b10111100110] = 16'b0000011111010011;
	exp_table[11'b10111100111] = 16'b0000011111011011;
	exp_table[11'b10111101000] = 16'b0000011111100010;
	exp_table[11'b10111101001] = 16'b0000011111101010;
	exp_table[11'b10111101010] = 16'b0000011111110010;
	exp_table[11'b10111101011] = 16'b0000011111111010;
	exp_table[11'b10111101100] = 16'b0000100000000010;
	exp_table[11'b10111101101] = 16'b0000100000001010;
	exp_table[11'b10111101110] = 16'b0000100000010010;
	exp_table[11'b10111101111] = 16'b0000100000011010;
	exp_table[11'b10111110000] = 16'b0000100000100010;
	exp_table[11'b10111110001] = 16'b0000100000101011;
	exp_table[11'b10111110010] = 16'b0000100000110011;
	exp_table[11'b10111110011] = 16'b0000100000111011;
	exp_table[11'b10111110100] = 16'b0000100001000011;
	exp_table[11'b10111110101] = 16'b0000100001001100;
	exp_table[11'b10111110110] = 16'b0000100001010100;
	exp_table[11'b10111110111] = 16'b0000100001011100;
	exp_table[11'b10111111000] = 16'b0000100001100101;
	exp_table[11'b10111111001] = 16'b0000100001101101;
	exp_table[11'b10111111010] = 16'b0000100001110101;
	exp_table[11'b10111111011] = 16'b0000100001111110;
	exp_table[11'b10111111100] = 16'b0000100010000110;
	exp_table[11'b10111111101] = 16'b0000100010001111;
	exp_table[11'b10111111110] = 16'b0000100010011000;
	exp_table[11'b10111111111] = 16'b0000100010100000;
	exp_table[11'b11000000000] = 16'b0000100010101001;
	exp_table[11'b11000000001] = 16'b0000100010110010;
	exp_table[11'b11000000010] = 16'b0000100010111010;
	exp_table[11'b11000000011] = 16'b0000100011000011;
	exp_table[11'b11000000100] = 16'b0000100011001100;
	exp_table[11'b11000000101] = 16'b0000100011010101;
	exp_table[11'b11000000110] = 16'b0000100011011101;
	exp_table[11'b11000000111] = 16'b0000100011100110;
	exp_table[11'b11000001000] = 16'b0000100011101111;
	exp_table[11'b11000001001] = 16'b0000100011111000;
	exp_table[11'b11000001010] = 16'b0000100100000001;
	exp_table[11'b11000001011] = 16'b0000100100001010;
	exp_table[11'b11000001100] = 16'b0000100100010011;
	exp_table[11'b11000001101] = 16'b0000100100011100;
	exp_table[11'b11000001110] = 16'b0000100100100101;
	exp_table[11'b11000001111] = 16'b0000100100101111;
	exp_table[11'b11000010000] = 16'b0000100100111000;
	exp_table[11'b11000010001] = 16'b0000100101000001;
	exp_table[11'b11000010010] = 16'b0000100101001010;
	exp_table[11'b11000010011] = 16'b0000100101010100;
	exp_table[11'b11000010100] = 16'b0000100101011101;
	exp_table[11'b11000010101] = 16'b0000100101100110;
	exp_table[11'b11000010110] = 16'b0000100101110000;
	exp_table[11'b11000010111] = 16'b0000100101111001;
	exp_table[11'b11000011000] = 16'b0000100110000011;
	exp_table[11'b11000011001] = 16'b0000100110001100;
	exp_table[11'b11000011010] = 16'b0000100110010110;
	exp_table[11'b11000011011] = 16'b0000100110011111;
	exp_table[11'b11000011100] = 16'b0000100110101001;
	exp_table[11'b11000011101] = 16'b0000100110110011;
	exp_table[11'b11000011110] = 16'b0000100110111101;
	exp_table[11'b11000011111] = 16'b0000100111000110;
	exp_table[11'b11000100000] = 16'b0000100111010000;
	exp_table[11'b11000100001] = 16'b0000100111011010;
	exp_table[11'b11000100010] = 16'b0000100111100100;
	exp_table[11'b11000100011] = 16'b0000100111101110;
	exp_table[11'b11000100100] = 16'b0000100111111000;
	exp_table[11'b11000100101] = 16'b0000101000000010;
	exp_table[11'b11000100110] = 16'b0000101000001100;
	exp_table[11'b11000100111] = 16'b0000101000010110;
	exp_table[11'b11000101000] = 16'b0000101000100000;
	exp_table[11'b11000101001] = 16'b0000101000101010;
	exp_table[11'b11000101010] = 16'b0000101000110100;
	exp_table[11'b11000101011] = 16'b0000101000111110;
	exp_table[11'b11000101100] = 16'b0000101001001001;
	exp_table[11'b11000101101] = 16'b0000101001010011;
	exp_table[11'b11000101110] = 16'b0000101001011101;
	exp_table[11'b11000101111] = 16'b0000101001101000;
	exp_table[11'b11000110000] = 16'b0000101001110010;
	exp_table[11'b11000110001] = 16'b0000101001111101;
	exp_table[11'b11000110010] = 16'b0000101010000111;
	exp_table[11'b11000110011] = 16'b0000101010010010;
	exp_table[11'b11000110100] = 16'b0000101010011100;
	exp_table[11'b11000110101] = 16'b0000101010100111;
	exp_table[11'b11000110110] = 16'b0000101010110010;
	exp_table[11'b11000110111] = 16'b0000101010111100;
	exp_table[11'b11000111000] = 16'b0000101011000111;
	exp_table[11'b11000111001] = 16'b0000101011010010;
	exp_table[11'b11000111010] = 16'b0000101011011101;
	exp_table[11'b11000111011] = 16'b0000101011101000;
	exp_table[11'b11000111100] = 16'b0000101011110010;
	exp_table[11'b11000111101] = 16'b0000101011111101;
	exp_table[11'b11000111110] = 16'b0000101100001000;
	exp_table[11'b11000111111] = 16'b0000101100010100;
	exp_table[11'b11001000000] = 16'b0000101100011111;
	exp_table[11'b11001000001] = 16'b0000101100101010;
	exp_table[11'b11001000010] = 16'b0000101100110101;
	exp_table[11'b11001000011] = 16'b0000101101000000;
	exp_table[11'b11001000100] = 16'b0000101101001011;
	exp_table[11'b11001000101] = 16'b0000101101010111;
	exp_table[11'b11001000110] = 16'b0000101101100010;
	exp_table[11'b11001000111] = 16'b0000101101101110;
	exp_table[11'b11001001000] = 16'b0000101101111001;
	exp_table[11'b11001001001] = 16'b0000101110000100;
	exp_table[11'b11001001010] = 16'b0000101110010000;
	exp_table[11'b11001001011] = 16'b0000101110011100;
	exp_table[11'b11001001100] = 16'b0000101110100111;
	exp_table[11'b11001001101] = 16'b0000101110110011;
	exp_table[11'b11001001110] = 16'b0000101110111111;
	exp_table[11'b11001001111] = 16'b0000101111001010;
	exp_table[11'b11001010000] = 16'b0000101111010110;
	exp_table[11'b11001010001] = 16'b0000101111100010;
	exp_table[11'b11001010010] = 16'b0000101111101110;
	exp_table[11'b11001010011] = 16'b0000101111111010;
	exp_table[11'b11001010100] = 16'b0000110000000110;
	exp_table[11'b11001010101] = 16'b0000110000010010;
	exp_table[11'b11001010110] = 16'b0000110000011110;
	exp_table[11'b11001010111] = 16'b0000110000101010;
	exp_table[11'b11001011000] = 16'b0000110000110110;
	exp_table[11'b11001011001] = 16'b0000110001000011;
	exp_table[11'b11001011010] = 16'b0000110001001111;
	exp_table[11'b11001011011] = 16'b0000110001011011;
	exp_table[11'b11001011100] = 16'b0000110001101000;
	exp_table[11'b11001011101] = 16'b0000110001110100;
	exp_table[11'b11001011110] = 16'b0000110010000001;
	exp_table[11'b11001011111] = 16'b0000110010001101;
	exp_table[11'b11001100000] = 16'b0000110010011010;
	exp_table[11'b11001100001] = 16'b0000110010100110;
	exp_table[11'b11001100010] = 16'b0000110010110011;
	exp_table[11'b11001100011] = 16'b0000110011000000;
	exp_table[11'b11001100100] = 16'b0000110011001101;
	exp_table[11'b11001100101] = 16'b0000110011011001;
	exp_table[11'b11001100110] = 16'b0000110011100110;
	exp_table[11'b11001100111] = 16'b0000110011110011;
	exp_table[11'b11001101000] = 16'b0000110100000000;
	exp_table[11'b11001101001] = 16'b0000110100001101;
	exp_table[11'b11001101010] = 16'b0000110100011010;
	exp_table[11'b11001101011] = 16'b0000110100100111;
	exp_table[11'b11001101100] = 16'b0000110100110101;
	exp_table[11'b11001101101] = 16'b0000110101000010;
	exp_table[11'b11001101110] = 16'b0000110101001111;
	exp_table[11'b11001101111] = 16'b0000110101011100;
	exp_table[11'b11001110000] = 16'b0000110101101010;
	exp_table[11'b11001110001] = 16'b0000110101110111;
	exp_table[11'b11001110010] = 16'b0000110110000101;
	exp_table[11'b11001110011] = 16'b0000110110010010;
	exp_table[11'b11001110100] = 16'b0000110110100000;
	exp_table[11'b11001110101] = 16'b0000110110101110;
	exp_table[11'b11001110110] = 16'b0000110110111011;
	exp_table[11'b11001110111] = 16'b0000110111001001;
	exp_table[11'b11001111000] = 16'b0000110111010111;
	exp_table[11'b11001111001] = 16'b0000110111100101;
	exp_table[11'b11001111010] = 16'b0000110111110011;
	exp_table[11'b11001111011] = 16'b0000111000000001;
	exp_table[11'b11001111100] = 16'b0000111000001111;
	exp_table[11'b11001111101] = 16'b0000111000011101;
	exp_table[11'b11001111110] = 16'b0000111000101011;
	exp_table[11'b11001111111] = 16'b0000111000111001;
	exp_table[11'b11010000000] = 16'b0000111001000111;
	exp_table[11'b11010000001] = 16'b0000111001010110;
	exp_table[11'b11010000010] = 16'b0000111001100100;
	exp_table[11'b11010000011] = 16'b0000111001110010;
	exp_table[11'b11010000100] = 16'b0000111010000001;
	exp_table[11'b11010000101] = 16'b0000111010001111;
	exp_table[11'b11010000110] = 16'b0000111010011110;
	exp_table[11'b11010000111] = 16'b0000111010101101;
	exp_table[11'b11010001000] = 16'b0000111010111011;
	exp_table[11'b11010001001] = 16'b0000111011001010;
	exp_table[11'b11010001010] = 16'b0000111011011001;
	exp_table[11'b11010001011] = 16'b0000111011101000;
	exp_table[11'b11010001100] = 16'b0000111011110111;
	exp_table[11'b11010001101] = 16'b0000111100000110;
	exp_table[11'b11010001110] = 16'b0000111100010101;
	exp_table[11'b11010001111] = 16'b0000111100100100;
	exp_table[11'b11010010000] = 16'b0000111100110011;
	exp_table[11'b11010010001] = 16'b0000111101000010;
	exp_table[11'b11010010010] = 16'b0000111101010010;
	exp_table[11'b11010010011] = 16'b0000111101100001;
	exp_table[11'b11010010100] = 16'b0000111101110000;
	exp_table[11'b11010010101] = 16'b0000111110000000;
	exp_table[11'b11010010110] = 16'b0000111110001111;
	exp_table[11'b11010010111] = 16'b0000111110011111;
	exp_table[11'b11010011000] = 16'b0000111110101111;
	exp_table[11'b11010011001] = 16'b0000111110111110;
	exp_table[11'b11010011010] = 16'b0000111111001110;
	exp_table[11'b11010011011] = 16'b0000111111011110;
	exp_table[11'b11010011100] = 16'b0000111111101110;
	exp_table[11'b11010011101] = 16'b0000111111111110;
	exp_table[11'b11010011110] = 16'b0001000000001110;
	exp_table[11'b11010011111] = 16'b0001000000011110;
	exp_table[11'b11010100000] = 16'b0001000000101110;
	exp_table[11'b11010100001] = 16'b0001000000111110;
	exp_table[11'b11010100010] = 16'b0001000001001111;
	exp_table[11'b11010100011] = 16'b0001000001011111;
	exp_table[11'b11010100100] = 16'b0001000001101111;
	exp_table[11'b11010100101] = 16'b0001000010000000;
	exp_table[11'b11010100110] = 16'b0001000010010000;
	exp_table[11'b11010100111] = 16'b0001000010100001;
	exp_table[11'b11010101000] = 16'b0001000010110010;
	exp_table[11'b11010101001] = 16'b0001000011000010;
	exp_table[11'b11010101010] = 16'b0001000011010011;
	exp_table[11'b11010101011] = 16'b0001000011100100;
	exp_table[11'b11010101100] = 16'b0001000011110101;
	exp_table[11'b11010101101] = 16'b0001000100000110;
	exp_table[11'b11010101110] = 16'b0001000100010111;
	exp_table[11'b11010101111] = 16'b0001000100101000;
	exp_table[11'b11010110000] = 16'b0001000100111001;
	exp_table[11'b11010110001] = 16'b0001000101001010;
	exp_table[11'b11010110010] = 16'b0001000101011100;
	exp_table[11'b11010110011] = 16'b0001000101101101;
	exp_table[11'b11010110100] = 16'b0001000101111111;
	exp_table[11'b11010110101] = 16'b0001000110010000;
	exp_table[11'b11010110110] = 16'b0001000110100010;
	exp_table[11'b11010110111] = 16'b0001000110110011;
	exp_table[11'b11010111000] = 16'b0001000111000101;
	exp_table[11'b11010111001] = 16'b0001000111010111;
	exp_table[11'b11010111010] = 16'b0001000111101001;
	exp_table[11'b11010111011] = 16'b0001000111111011;
	exp_table[11'b11010111100] = 16'b0001001000001101;
	exp_table[11'b11010111101] = 16'b0001001000011111;
	exp_table[11'b11010111110] = 16'b0001001000110001;
	exp_table[11'b11010111111] = 16'b0001001001000011;
	exp_table[11'b11011000000] = 16'b0001001001010110;
	exp_table[11'b11011000001] = 16'b0001001001101000;
	exp_table[11'b11011000010] = 16'b0001001001111010;
	exp_table[11'b11011000011] = 16'b0001001010001101;
	exp_table[11'b11011000100] = 16'b0001001010100000;
	exp_table[11'b11011000101] = 16'b0001001010110010;
	exp_table[11'b11011000110] = 16'b0001001011000101;
	exp_table[11'b11011000111] = 16'b0001001011011000;
	exp_table[11'b11011001000] = 16'b0001001011101011;
	exp_table[11'b11011001001] = 16'b0001001011111110;
	exp_table[11'b11011001010] = 16'b0001001100010001;
	exp_table[11'b11011001011] = 16'b0001001100100100;
	exp_table[11'b11011001100] = 16'b0001001100110111;
	exp_table[11'b11011001101] = 16'b0001001101001010;
	exp_table[11'b11011001110] = 16'b0001001101011101;
	exp_table[11'b11011001111] = 16'b0001001101110001;
	exp_table[11'b11011010000] = 16'b0001001110000100;
	exp_table[11'b11011010001] = 16'b0001001110011000;
	exp_table[11'b11011010010] = 16'b0001001110101100;
	exp_table[11'b11011010011] = 16'b0001001110111111;
	exp_table[11'b11011010100] = 16'b0001001111010011;
	exp_table[11'b11011010101] = 16'b0001001111100111;
	exp_table[11'b11011010110] = 16'b0001001111111011;
	exp_table[11'b11011010111] = 16'b0001010000001111;
	exp_table[11'b11011011000] = 16'b0001010000100011;
	exp_table[11'b11011011001] = 16'b0001010000110111;
	exp_table[11'b11011011010] = 16'b0001010001001011;
	exp_table[11'b11011011011] = 16'b0001010001100000;
	exp_table[11'b11011011100] = 16'b0001010001110100;
	exp_table[11'b11011011101] = 16'b0001010010001001;
	exp_table[11'b11011011110] = 16'b0001010010011101;
	exp_table[11'b11011011111] = 16'b0001010010110010;
	exp_table[11'b11011100000] = 16'b0001010011000111;
	exp_table[11'b11011100001] = 16'b0001010011011011;
	exp_table[11'b11011100010] = 16'b0001010011110000;
	exp_table[11'b11011100011] = 16'b0001010100000101;
	exp_table[11'b11011100100] = 16'b0001010100011010;
	exp_table[11'b11011100101] = 16'b0001010100110000;
	exp_table[11'b11011100110] = 16'b0001010101000101;
	exp_table[11'b11011100111] = 16'b0001010101011010;
	exp_table[11'b11011101000] = 16'b0001010101101111;
	exp_table[11'b11011101001] = 16'b0001010110000101;
	exp_table[11'b11011101010] = 16'b0001010110011010;
	exp_table[11'b11011101011] = 16'b0001010110110000;
	exp_table[11'b11011101100] = 16'b0001010111000110;
	exp_table[11'b11011101101] = 16'b0001010111011100;
	exp_table[11'b11011101110] = 16'b0001010111110010;
	exp_table[11'b11011101111] = 16'b0001011000001000;
	exp_table[11'b11011110000] = 16'b0001011000011110;
	exp_table[11'b11011110001] = 16'b0001011000110100;
	exp_table[11'b11011110010] = 16'b0001011001001010;
	exp_table[11'b11011110011] = 16'b0001011001100000;
	exp_table[11'b11011110100] = 16'b0001011001110111;
	exp_table[11'b11011110101] = 16'b0001011010001101;
	exp_table[11'b11011110110] = 16'b0001011010100100;
	exp_table[11'b11011110111] = 16'b0001011010111011;
	exp_table[11'b11011111000] = 16'b0001011011010001;
	exp_table[11'b11011111001] = 16'b0001011011101000;
	exp_table[11'b11011111010] = 16'b0001011011111111;
	exp_table[11'b11011111011] = 16'b0001011100010110;
	exp_table[11'b11011111100] = 16'b0001011100101101;
	exp_table[11'b11011111101] = 16'b0001011101000101;
	exp_table[11'b11011111110] = 16'b0001011101011100;
	exp_table[11'b11011111111] = 16'b0001011101110011;
	exp_table[11'b11100000000] = 16'b0001011110001011;
	exp_table[11'b11100000001] = 16'b0001011110100010;
	exp_table[11'b11100000010] = 16'b0001011110111010;
	exp_table[11'b11100000011] = 16'b0001011111010010;
	exp_table[11'b11100000100] = 16'b0001011111101010;
	exp_table[11'b11100000101] = 16'b0001100000000010;
	exp_table[11'b11100000110] = 16'b0001100000011010;
	exp_table[11'b11100000111] = 16'b0001100000110010;
	exp_table[11'b11100001000] = 16'b0001100001001010;
	exp_table[11'b11100001001] = 16'b0001100001100011;
	exp_table[11'b11100001010] = 16'b0001100001111011;
	exp_table[11'b11100001011] = 16'b0001100010010011;
	exp_table[11'b11100001100] = 16'b0001100010101100;
	exp_table[11'b11100001101] = 16'b0001100011000101;
	exp_table[11'b11100001110] = 16'b0001100011011110;
	exp_table[11'b11100001111] = 16'b0001100011110111;
	exp_table[11'b11100010000] = 16'b0001100100010000;
	exp_table[11'b11100010001] = 16'b0001100100101001;
	exp_table[11'b11100010010] = 16'b0001100101000010;
	exp_table[11'b11100010011] = 16'b0001100101011011;
	exp_table[11'b11100010100] = 16'b0001100101110101;
	exp_table[11'b11100010101] = 16'b0001100110001110;
	exp_table[11'b11100010110] = 16'b0001100110101000;
	exp_table[11'b11100010111] = 16'b0001100111000001;
	exp_table[11'b11100011000] = 16'b0001100111011011;
	exp_table[11'b11100011001] = 16'b0001100111110101;
	exp_table[11'b11100011010] = 16'b0001101000001111;
	exp_table[11'b11100011011] = 16'b0001101000101001;
	exp_table[11'b11100011100] = 16'b0001101001000011;
	exp_table[11'b11100011101] = 16'b0001101001011110;
	exp_table[11'b11100011110] = 16'b0001101001111000;
	exp_table[11'b11100011111] = 16'b0001101010010011;
	exp_table[11'b11100100000] = 16'b0001101010101101;
	exp_table[11'b11100100001] = 16'b0001101011001000;
	exp_table[11'b11100100010] = 16'b0001101011100011;
	exp_table[11'b11100100011] = 16'b0001101011111110;
	exp_table[11'b11100100100] = 16'b0001101100011001;
	exp_table[11'b11100100101] = 16'b0001101100110100;
	exp_table[11'b11100100110] = 16'b0001101101001111;
	exp_table[11'b11100100111] = 16'b0001101101101011;
	exp_table[11'b11100101000] = 16'b0001101110000110;
	exp_table[11'b11100101001] = 16'b0001101110100010;
	exp_table[11'b11100101010] = 16'b0001101110111101;
	exp_table[11'b11100101011] = 16'b0001101111011001;
	exp_table[11'b11100101100] = 16'b0001101111110101;
	exp_table[11'b11100101101] = 16'b0001110000010001;
	exp_table[11'b11100101110] = 16'b0001110000101101;
	exp_table[11'b11100101111] = 16'b0001110001001010;
	exp_table[11'b11100110000] = 16'b0001110001100110;
	exp_table[11'b11100110001] = 16'b0001110010000010;
	exp_table[11'b11100110010] = 16'b0001110010011111;
	exp_table[11'b11100110011] = 16'b0001110010111100;
	exp_table[11'b11100110100] = 16'b0001110011011000;
	exp_table[11'b11100110101] = 16'b0001110011110101;
	exp_table[11'b11100110110] = 16'b0001110100010010;
	exp_table[11'b11100110111] = 16'b0001110100101111;
	exp_table[11'b11100111000] = 16'b0001110101001101;
	exp_table[11'b11100111001] = 16'b0001110101101010;
	exp_table[11'b11100111010] = 16'b0001110110000111;
	exp_table[11'b11100111011] = 16'b0001110110100101;
	exp_table[11'b11100111100] = 16'b0001110111000011;
	exp_table[11'b11100111101] = 16'b0001110111100001;
	exp_table[11'b11100111110] = 16'b0001110111111111;
	exp_table[11'b11100111111] = 16'b0001111000011101;
	exp_table[11'b11101000000] = 16'b0001111000111011;
	exp_table[11'b11101000001] = 16'b0001111001011001;
	exp_table[11'b11101000010] = 16'b0001111001110111;
	exp_table[11'b11101000011] = 16'b0001111010010110;
	exp_table[11'b11101000100] = 16'b0001111010110101;
	exp_table[11'b11101000101] = 16'b0001111011010011;
	exp_table[11'b11101000110] = 16'b0001111011110010;
	exp_table[11'b11101000111] = 16'b0001111100010001;
	exp_table[11'b11101001000] = 16'b0001111100110000;
	exp_table[11'b11101001001] = 16'b0001111101010000;
	exp_table[11'b11101001010] = 16'b0001111101101111;
	exp_table[11'b11101001011] = 16'b0001111110001111;
	exp_table[11'b11101001100] = 16'b0001111110101110;
	exp_table[11'b11101001101] = 16'b0001111111001110;
	exp_table[11'b11101001110] = 16'b0001111111101110;
	exp_table[11'b11101001111] = 16'b0010000000001110;
	exp_table[11'b11101010000] = 16'b0010000000101110;
	exp_table[11'b11101010001] = 16'b0010000001001110;
	exp_table[11'b11101010010] = 16'b0010000001101111;
	exp_table[11'b11101010011] = 16'b0010000010001111;
	exp_table[11'b11101010100] = 16'b0010000010110000;
	exp_table[11'b11101010101] = 16'b0010000011010000;
	exp_table[11'b11101010110] = 16'b0010000011110001;
	exp_table[11'b11101010111] = 16'b0010000100010010;
	exp_table[11'b11101011000] = 16'b0010000100110011;
	exp_table[11'b11101011001] = 16'b0010000101010101;
	exp_table[11'b11101011010] = 16'b0010000101110110;
	exp_table[11'b11101011011] = 16'b0010000110011000;
	exp_table[11'b11101011100] = 16'b0010000110111001;
	exp_table[11'b11101011101] = 16'b0010000111011011;
	exp_table[11'b11101011110] = 16'b0010000111111101;
	exp_table[11'b11101011111] = 16'b0010001000011111;
	exp_table[11'b11101100000] = 16'b0010001001000001;
	exp_table[11'b11101100001] = 16'b0010001001100100;
	exp_table[11'b11101100010] = 16'b0010001010000110;
	exp_table[11'b11101100011] = 16'b0010001010101001;
	exp_table[11'b11101100100] = 16'b0010001011001011;
	exp_table[11'b11101100101] = 16'b0010001011101110;
	exp_table[11'b11101100110] = 16'b0010001100010001;
	exp_table[11'b11101100111] = 16'b0010001100110100;
	exp_table[11'b11101101000] = 16'b0010001101011000;
	exp_table[11'b11101101001] = 16'b0010001101111011;
	exp_table[11'b11101101010] = 16'b0010001110011111;
	exp_table[11'b11101101011] = 16'b0010001111000010;
	exp_table[11'b11101101100] = 16'b0010001111100110;
	exp_table[11'b11101101101] = 16'b0010010000001010;
	exp_table[11'b11101101110] = 16'b0010010000101110;
	exp_table[11'b11101101111] = 16'b0010010001010010;
	exp_table[11'b11101110000] = 16'b0010010001110111;
	exp_table[11'b11101110001] = 16'b0010010010011011;
	exp_table[11'b11101110010] = 16'b0010010011000000;
	exp_table[11'b11101110011] = 16'b0010010011100101;
	exp_table[11'b11101110100] = 16'b0010010100001010;
	exp_table[11'b11101110101] = 16'b0010010100101111;
	exp_table[11'b11101110110] = 16'b0010010101010100;
	exp_table[11'b11101110111] = 16'b0010010101111010;
	exp_table[11'b11101111000] = 16'b0010010110011111;
	exp_table[11'b11101111001] = 16'b0010010111000101;
	exp_table[11'b11101111010] = 16'b0010010111101011;
	exp_table[11'b11101111011] = 16'b0010011000010001;
	exp_table[11'b11101111100] = 16'b0010011000110111;
	exp_table[11'b11101111101] = 16'b0010011001011101;
	exp_table[11'b11101111110] = 16'b0010011010000100;
	exp_table[11'b11101111111] = 16'b0010011010101010;
	exp_table[11'b11110000000] = 16'b0010011011010001;
	exp_table[11'b11110000001] = 16'b0010011011111000;
	exp_table[11'b11110000010] = 16'b0010011100011111;
	exp_table[11'b11110000011] = 16'b0010011101000110;
	exp_table[11'b11110000100] = 16'b0010011101101101;
	exp_table[11'b11110000101] = 16'b0010011110010101;
	exp_table[11'b11110000110] = 16'b0010011110111101;
	exp_table[11'b11110000111] = 16'b0010011111100100;
	exp_table[11'b11110001000] = 16'b0010100000001100;
	exp_table[11'b11110001001] = 16'b0010100000110100;
	exp_table[11'b11110001010] = 16'b0010100001011101;
	exp_table[11'b11110001011] = 16'b0010100010000101;
	exp_table[11'b11110001100] = 16'b0010100010101110;
	exp_table[11'b11110001101] = 16'b0010100011010111;
	exp_table[11'b11110001110] = 16'b0010100011111111;
	exp_table[11'b11110001111] = 16'b0010100100101001;
	exp_table[11'b11110010000] = 16'b0010100101010010;
	exp_table[11'b11110010001] = 16'b0010100101111011;
	exp_table[11'b11110010010] = 16'b0010100110100101;
	exp_table[11'b11110010011] = 16'b0010100111001110;
	exp_table[11'b11110010100] = 16'b0010100111111000;
	exp_table[11'b11110010101] = 16'b0010101000100010;
	exp_table[11'b11110010110] = 16'b0010101001001101;
	exp_table[11'b11110010111] = 16'b0010101001110111;
	exp_table[11'b11110011000] = 16'b0010101010100010;
	exp_table[11'b11110011001] = 16'b0010101011001100;
	exp_table[11'b11110011010] = 16'b0010101011110111;
	exp_table[11'b11110011011] = 16'b0010101100100010;
	exp_table[11'b11110011100] = 16'b0010101101001101;
	exp_table[11'b11110011101] = 16'b0010101101111001;
	exp_table[11'b11110011110] = 16'b0010101110100100;
	exp_table[11'b11110011111] = 16'b0010101111010000;
	exp_table[11'b11110100000] = 16'b0010101111111100;
	exp_table[11'b11110100001] = 16'b0010110000101000;
	exp_table[11'b11110100010] = 16'b0010110001010100;
	exp_table[11'b11110100011] = 16'b0010110010000001;
	exp_table[11'b11110100100] = 16'b0010110010101101;
	exp_table[11'b11110100101] = 16'b0010110011011010;
	exp_table[11'b11110100110] = 16'b0010110100000111;
	exp_table[11'b11110100111] = 16'b0010110100110100;
	exp_table[11'b11110101000] = 16'b0010110101100001;
	exp_table[11'b11110101001] = 16'b0010110110001111;
	exp_table[11'b11110101010] = 16'b0010110110111101;
	exp_table[11'b11110101011] = 16'b0010110111101010;
	exp_table[11'b11110101100] = 16'b0010111000011000;
	exp_table[11'b11110101101] = 16'b0010111001000111;
	exp_table[11'b11110101110] = 16'b0010111001110101;
	exp_table[11'b11110101111] = 16'b0010111010100100;
	exp_table[11'b11110110000] = 16'b0010111011010010;
	exp_table[11'b11110110001] = 16'b0010111100000001;
	exp_table[11'b11110110010] = 16'b0010111100110000;
	exp_table[11'b11110110011] = 16'b0010111101100000;
	exp_table[11'b11110110100] = 16'b0010111110001111;
	exp_table[11'b11110110101] = 16'b0010111110111111;
	exp_table[11'b11110110110] = 16'b0010111111101111;
	exp_table[11'b11110110111] = 16'b0011000000011111;
	exp_table[11'b11110111000] = 16'b0011000001001111;
	exp_table[11'b11110111001] = 16'b0011000001111111;
	exp_table[11'b11110111010] = 16'b0011000010110000;
	exp_table[11'b11110111011] = 16'b0011000011100001;
	exp_table[11'b11110111100] = 16'b0011000100010010;
	exp_table[11'b11110111101] = 16'b0011000101000011;
	exp_table[11'b11110111110] = 16'b0011000101110100;
	exp_table[11'b11110111111] = 16'b0011000110100110;
	exp_table[11'b11111000000] = 16'b0011000111010111;
	exp_table[11'b11111000001] = 16'b0011001000001001;
	exp_table[11'b11111000010] = 16'b0011001000111011;
	exp_table[11'b11111000011] = 16'b0011001001101110;
	exp_table[11'b11111000100] = 16'b0011001010100000;
	exp_table[11'b11111000101] = 16'b0011001011010011;
	exp_table[11'b11111000110] = 16'b0011001100000110;
	exp_table[11'b11111000111] = 16'b0011001100111001;
	exp_table[11'b11111001000] = 16'b0011001101101100;
	exp_table[11'b11111001001] = 16'b0011001110100000;
	exp_table[11'b11111001010] = 16'b0011001111010100;
	exp_table[11'b11111001011] = 16'b0011010000001000;
	exp_table[11'b11111001100] = 16'b0011010000111100;
	exp_table[11'b11111001101] = 16'b0011010001110000;
	exp_table[11'b11111001110] = 16'b0011010010100101;
	exp_table[11'b11111001111] = 16'b0011010011011001;
	exp_table[11'b11111010000] = 16'b0011010100001110;
	exp_table[11'b11111010001] = 16'b0011010101000011;
	exp_table[11'b11111010010] = 16'b0011010101111001;
	exp_table[11'b11111010011] = 16'b0011010110101110;
	exp_table[11'b11111010100] = 16'b0011010111100100;
	exp_table[11'b11111010101] = 16'b0011011000011010;
	exp_table[11'b11111010110] = 16'b0011011001010000;
	exp_table[11'b11111010111] = 16'b0011011010000111;
	exp_table[11'b11111011000] = 16'b0011011010111101;
	exp_table[11'b11111011001] = 16'b0011011011110100;
	exp_table[11'b11111011010] = 16'b0011011100101011;
	exp_table[11'b11111011011] = 16'b0011011101100011;
	exp_table[11'b11111011100] = 16'b0011011110011010;
	exp_table[11'b11111011101] = 16'b0011011111010010;
	exp_table[11'b11111011110] = 16'b0011100000001010;
	exp_table[11'b11111011111] = 16'b0011100001000010;
	exp_table[11'b11111100000] = 16'b0011100001111010;
	exp_table[11'b11111100001] = 16'b0011100010110011;
	exp_table[11'b11111100010] = 16'b0011100011101100;
	exp_table[11'b11111100011] = 16'b0011100100100101;
	exp_table[11'b11111100100] = 16'b0011100101011110;
	exp_table[11'b11111100101] = 16'b0011100110011000;
	exp_table[11'b11111100110] = 16'b0011100111010001;
	exp_table[11'b11111100111] = 16'b0011101000001011;
	exp_table[11'b11111101000] = 16'b0011101001000101;
	exp_table[11'b11111101001] = 16'b0011101010000000;
	exp_table[11'b11111101010] = 16'b0011101010111010;
	exp_table[11'b11111101011] = 16'b0011101011110101;
	exp_table[11'b11111101100] = 16'b0011101100110000;
	exp_table[11'b11111101101] = 16'b0011101101101100;
	exp_table[11'b11111101110] = 16'b0011101110100111;
	exp_table[11'b11111101111] = 16'b0011101111100011;
	exp_table[11'b11111110000] = 16'b0011110000011111;
	exp_table[11'b11111110001] = 16'b0011110001011011;
	exp_table[11'b11111110010] = 16'b0011110010011000;
	exp_table[11'b11111110011] = 16'b0011110011010100;
	exp_table[11'b11111110100] = 16'b0011110100010001;
	exp_table[11'b11111110101] = 16'b0011110101001110;
	exp_table[11'b11111110110] = 16'b0011110110001100;
	exp_table[11'b11111110111] = 16'b0011110111001010;
	exp_table[11'b11111111000] = 16'b0011111000000111;
	exp_table[11'b11111111001] = 16'b0011111001000110;
	exp_table[11'b11111111010] = 16'b0011111010000100;
	exp_table[11'b11111111011] = 16'b0011111011000011;
	exp_table[11'b11111111100] = 16'b0011111100000001;
	exp_table[11'b11111111101] = 16'b0011111101000001;
	exp_table[11'b11111111110] = 16'b0011111110000000;
	exp_table[11'b11111111111] = 16'b0011111111000000;
	exp_table[11'b00000000000] = 16'b0100000000000000;
	exp_table[11'b00000000001] = 16'b0100000001000000;
	exp_table[11'b00000000010] = 16'b0100000010000000;
	exp_table[11'b00000000011] = 16'b0100000011000001;
	exp_table[11'b00000000100] = 16'b0100000100000010;
	exp_table[11'b00000000101] = 16'b0100000101000011;
	exp_table[11'b00000000110] = 16'b0100000110000100;
	exp_table[11'b00000000111] = 16'b0100000111000110;
	exp_table[11'b00000001000] = 16'b0100001000001000;
	exp_table[11'b00000001001] = 16'b0100001001001010;
	exp_table[11'b00000001010] = 16'b0100001010001100;
	exp_table[11'b00000001011] = 16'b0100001011001111;
	exp_table[11'b00000001100] = 16'b0100001100010010;
	exp_table[11'b00000001101] = 16'b0100001101010101;
	exp_table[11'b00000001110] = 16'b0100001110011000;
	exp_table[11'b00000001111] = 16'b0100001111011100;
	exp_table[11'b00000010000] = 16'b0100010000100000;
	exp_table[11'b00000010001] = 16'b0100010001100100;
	exp_table[11'b00000010010] = 16'b0100010010101001;
	exp_table[11'b00000010011] = 16'b0100010011101110;
	exp_table[11'b00000010100] = 16'b0100010100110011;
	exp_table[11'b00000010101] = 16'b0100010101111000;
	exp_table[11'b00000010110] = 16'b0100010110111110;
	exp_table[11'b00000010111] = 16'b0100011000000100;
	exp_table[11'b00000011000] = 16'b0100011001001010;
	exp_table[11'b00000011001] = 16'b0100011010010000;
	exp_table[11'b00000011010] = 16'b0100011011010111;
	exp_table[11'b00000011011] = 16'b0100011100011110;
	exp_table[11'b00000011100] = 16'b0100011101100101;
	exp_table[11'b00000011101] = 16'b0100011110101101;
	exp_table[11'b00000011110] = 16'b0100011111110101;
	exp_table[11'b00000011111] = 16'b0100100000111101;
	exp_table[11'b00000100000] = 16'b0100100010000101;
	exp_table[11'b00000100001] = 16'b0100100011001110;
	exp_table[11'b00000100010] = 16'b0100100100010111;
	exp_table[11'b00000100011] = 16'b0100100101100000;
	exp_table[11'b00000100100] = 16'b0100100110101001;
	exp_table[11'b00000100101] = 16'b0100100111110011;
	exp_table[11'b00000100110] = 16'b0100101000111101;
	exp_table[11'b00000100111] = 16'b0100101010001000;
	exp_table[11'b00000101000] = 16'b0100101011010010;
	exp_table[11'b00000101001] = 16'b0100101100011101;
	exp_table[11'b00000101010] = 16'b0100101101101001;
	exp_table[11'b00000101011] = 16'b0100101110110100;
	exp_table[11'b00000101100] = 16'b0100110000000000;
	exp_table[11'b00000101101] = 16'b0100110001001100;
	exp_table[11'b00000101110] = 16'b0100110010011001;
	exp_table[11'b00000101111] = 16'b0100110011100101;
	exp_table[11'b00000110000] = 16'b0100110100110010;
	exp_table[11'b00000110001] = 16'b0100110110000000;
	exp_table[11'b00000110010] = 16'b0100110111001101;
	exp_table[11'b00000110011] = 16'b0100111000011011;
	exp_table[11'b00000110100] = 16'b0100111001101010;
	exp_table[11'b00000110101] = 16'b0100111010111000;
	exp_table[11'b00000110110] = 16'b0100111100000111;
	exp_table[11'b00000110111] = 16'b0100111101010110;
	exp_table[11'b00000111000] = 16'b0100111110100110;
	exp_table[11'b00000111001] = 16'b0100111111110110;
	exp_table[11'b00000111010] = 16'b0101000001000110;
	exp_table[11'b00000111011] = 16'b0101000010010110;
	exp_table[11'b00000111100] = 16'b0101000011100111;
	exp_table[11'b00000111101] = 16'b0101000100111000;
	exp_table[11'b00000111110] = 16'b0101000110001001;
	exp_table[11'b00000111111] = 16'b0101000111011011;
	exp_table[11'b00001000000] = 16'b0101001000101101;
	exp_table[11'b00001000001] = 16'b0101001001111111;
	exp_table[11'b00001000010] = 16'b0101001011010010;
	exp_table[11'b00001000011] = 16'b0101001100100101;
	exp_table[11'b00001000100] = 16'b0101001101111000;
	exp_table[11'b00001000101] = 16'b0101001111001100;
	exp_table[11'b00001000110] = 16'b0101010000100000;
	exp_table[11'b00001000111] = 16'b0101010001110100;
	exp_table[11'b00001001000] = 16'b0101010011001001;
	exp_table[11'b00001001001] = 16'b0101010100011110;
	exp_table[11'b00001001010] = 16'b0101010101110011;
	exp_table[11'b00001001011] = 16'b0101010111001001;
	exp_table[11'b00001001100] = 16'b0101011000011111;
	exp_table[11'b00001001101] = 16'b0101011001110101;
	exp_table[11'b00001001110] = 16'b0101011011001011;
	exp_table[11'b00001001111] = 16'b0101011100100010;
	exp_table[11'b00001010000] = 16'b0101011101111010;
	exp_table[11'b00001010001] = 16'b0101011111010001;
	exp_table[11'b00001010010] = 16'b0101100000101001;
	exp_table[11'b00001010011] = 16'b0101100010000010;
	exp_table[11'b00001010100] = 16'b0101100011011010;
	exp_table[11'b00001010101] = 16'b0101100100110011;
	exp_table[11'b00001010110] = 16'b0101100110001101;
	exp_table[11'b00001010111] = 16'b0101100111100111;
	exp_table[11'b00001011000] = 16'b0101101001000001;
	exp_table[11'b00001011001] = 16'b0101101010011011;
	exp_table[11'b00001011010] = 16'b0101101011110110;
	exp_table[11'b00001011011] = 16'b0101101101010001;
	exp_table[11'b00001011100] = 16'b0101101110101100;
	exp_table[11'b00001011101] = 16'b0101110000001000;
	exp_table[11'b00001011110] = 16'b0101110001100101;
	exp_table[11'b00001011111] = 16'b0101110011000001;
	exp_table[11'b00001100000] = 16'b0101110100011110;
	exp_table[11'b00001100001] = 16'b0101110101111011;
	exp_table[11'b00001100010] = 16'b0101110111011001;
	exp_table[11'b00001100011] = 16'b0101111000110111;
	exp_table[11'b00001100100] = 16'b0101111010010101;
	exp_table[11'b00001100101] = 16'b0101111011110100;
	exp_table[11'b00001100110] = 16'b0101111101010011;
	exp_table[11'b00001100111] = 16'b0101111110110011;
	exp_table[11'b00001101000] = 16'b0110000000010011;
	exp_table[11'b00001101001] = 16'b0110000001110011;
	exp_table[11'b00001101010] = 16'b0110000011010100;
	exp_table[11'b00001101011] = 16'b0110000100110101;
	exp_table[11'b00001101100] = 16'b0110000110010110;
	exp_table[11'b00001101101] = 16'b0110000111111000;
	exp_table[11'b00001101110] = 16'b0110001001011010;
	exp_table[11'b00001101111] = 16'b0110001010111101;
	exp_table[11'b00001110000] = 16'b0110001100100000;
	exp_table[11'b00001110001] = 16'b0110001110000011;
	exp_table[11'b00001110010] = 16'b0110001111100111;
	exp_table[11'b00001110011] = 16'b0110010001001011;
	exp_table[11'b00001110100] = 16'b0110010010101111;
	exp_table[11'b00001110101] = 16'b0110010100010100;
	exp_table[11'b00001110110] = 16'b0110010101111001;
	exp_table[11'b00001110111] = 16'b0110010111011111;
	exp_table[11'b00001111000] = 16'b0110011001000101;
	exp_table[11'b00001111001] = 16'b0110011010101100;
	exp_table[11'b00001111010] = 16'b0110011100010010;
	exp_table[11'b00001111011] = 16'b0110011101111010;
	exp_table[11'b00001111100] = 16'b0110011111100001;
	exp_table[11'b00001111101] = 16'b0110100001001001;
	exp_table[11'b00001111110] = 16'b0110100010110010;
	exp_table[11'b00001111111] = 16'b0110100100011011;
	exp_table[11'b00010000000] = 16'b0110100110000100;
	exp_table[11'b00010000001] = 16'b0110100111101110;
	exp_table[11'b00010000010] = 16'b0110101001011000;
	exp_table[11'b00010000011] = 16'b0110101011000011;
	exp_table[11'b00010000100] = 16'b0110101100101110;
	exp_table[11'b00010000101] = 16'b0110101110011001;
	exp_table[11'b00010000110] = 16'b0110110000000101;
	exp_table[11'b00010000111] = 16'b0110110001110001;
	exp_table[11'b00010001000] = 16'b0110110011011110;
	exp_table[11'b00010001001] = 16'b0110110101001011;
	exp_table[11'b00010001010] = 16'b0110110110111000;
	exp_table[11'b00010001011] = 16'b0110111000100110;
	exp_table[11'b00010001100] = 16'b0110111010010101;
	exp_table[11'b00010001101] = 16'b0110111100000011;
	exp_table[11'b00010001110] = 16'b0110111101110011;
	exp_table[11'b00010001111] = 16'b0110111111100010;
	exp_table[11'b00010010000] = 16'b0111000001010010;
	exp_table[11'b00010010001] = 16'b0111000011000011;
	exp_table[11'b00010010010] = 16'b0111000100110100;
	exp_table[11'b00010010011] = 16'b0111000110100101;
	exp_table[11'b00010010100] = 16'b0111001000010111;
	exp_table[11'b00010010101] = 16'b0111001010001001;
	exp_table[11'b00010010110] = 16'b0111001011111100;
	exp_table[11'b00010010111] = 16'b0111001101101111;
	exp_table[11'b00010011000] = 16'b0111001111100011;
	exp_table[11'b00010011001] = 16'b0111010001010111;
	exp_table[11'b00010011010] = 16'b0111010011001100;
	exp_table[11'b00010011011] = 16'b0111010101000001;
	exp_table[11'b00010011100] = 16'b0111010110110110;
	exp_table[11'b00010011101] = 16'b0111011000101100;
	exp_table[11'b00010011110] = 16'b0111011010100011;
	exp_table[11'b00010011111] = 16'b0111011100011010;
	exp_table[11'b00010100000] = 16'b0111011110010001;
	exp_table[11'b00010100001] = 16'b0111100000001001;
	exp_table[11'b00010100010] = 16'b0111100010000001;
	exp_table[11'b00010100011] = 16'b0111100011111010;
	exp_table[11'b00010100100] = 16'b0111100101110011;
	exp_table[11'b00010100101] = 16'b0111100111101101;
	exp_table[11'b00010100110] = 16'b0111101001100111;
	exp_table[11'b00010100111] = 16'b0111101011100001;
	exp_table[11'b00010101000] = 16'b0111101101011100;
	exp_table[11'b00010101001] = 16'b0111101111011000;
	exp_table[11'b00010101010] = 16'b0111110001010100;
	exp_table[11'b00010101011] = 16'b0111110011010001;
	exp_table[11'b00010101100] = 16'b0111110101001110;
	exp_table[11'b00010101101] = 16'b0111110111001011;
	exp_table[11'b00010101110] = 16'b0111111001001001;
	exp_table[11'b00010101111] = 16'b0111111011001000;
	exp_table[11'b00010110000] = 16'b0111111101000111;
	exp_table[11'b00010110001] = 16'b0111111111000111;
	exp_table[11'b00010110010] = 16'b1000000001000111;
	exp_table[11'b00010110011] = 16'b1000000011000111;
	exp_table[11'b00010110100] = 16'b1000000101001000;
	exp_table[11'b00010110101] = 16'b1000000111001010;
	exp_table[11'b00010110110] = 16'b1000001001001100;
	exp_table[11'b00010110111] = 16'b1000001011001110;
	exp_table[11'b00010111000] = 16'b1000001101010001;
	exp_table[11'b00010111001] = 16'b1000001111010101;
	exp_table[11'b00010111010] = 16'b1000010001011001;
	exp_table[11'b00010111011] = 16'b1000010011011110;
	exp_table[11'b00010111100] = 16'b1000010101100011;
	exp_table[11'b00010111101] = 16'b1000010111101000;
	exp_table[11'b00010111110] = 16'b1000011001101111;
	exp_table[11'b00010111111] = 16'b1000011011110101;
	exp_table[11'b00011000000] = 16'b1000011101111100;
	exp_table[11'b00011000001] = 16'b1000100000000100;
	exp_table[11'b00011000010] = 16'b1000100010001100;
	exp_table[11'b00011000011] = 16'b1000100100010101;
	exp_table[11'b00011000100] = 16'b1000100110011111;
	exp_table[11'b00011000101] = 16'b1000101000101001;
	exp_table[11'b00011000110] = 16'b1000101010110011;
	exp_table[11'b00011000111] = 16'b1000101100111110;
	exp_table[11'b00011001000] = 16'b1000101111001001;
	exp_table[11'b00011001001] = 16'b1000110001010110;
	exp_table[11'b00011001010] = 16'b1000110011100010;
	exp_table[11'b00011001011] = 16'b1000110101101111;
	exp_table[11'b00011001100] = 16'b1000110111111101;
	exp_table[11'b00011001101] = 16'b1000111010001011;
	exp_table[11'b00011001110] = 16'b1000111100011010;
	exp_table[11'b00011001111] = 16'b1000111110101001;
	exp_table[11'b00011010000] = 16'b1001000000111001;
	exp_table[11'b00011010001] = 16'b1001000011001010;
	exp_table[11'b00011010010] = 16'b1001000101011011;
	exp_table[11'b00011010011] = 16'b1001000111101101;
	exp_table[11'b00011010100] = 16'b1001001001111111;
	exp_table[11'b00011010101] = 16'b1001001100010010;
	exp_table[11'b00011010110] = 16'b1001001110100101;
	exp_table[11'b00011010111] = 16'b1001010000111001;
	exp_table[11'b00011011000] = 16'b1001010011001101;
	exp_table[11'b00011011001] = 16'b1001010101100011;
	exp_table[11'b00011011010] = 16'b1001010111111000;
	exp_table[11'b00011011011] = 16'b1001011010001110;
	exp_table[11'b00011011100] = 16'b1001011100100101;
	exp_table[11'b00011011101] = 16'b1001011110111101;
	exp_table[11'b00011011110] = 16'b1001100001010101;
	exp_table[11'b00011011111] = 16'b1001100011101101;
	exp_table[11'b00011100000] = 16'b1001100110000111;
	exp_table[11'b00011100001] = 16'b1001101000100001;
	exp_table[11'b00011100010] = 16'b1001101010111011;
	exp_table[11'b00011100011] = 16'b1001101101010110;
	exp_table[11'b00011100100] = 16'b1001101111110010;
	exp_table[11'b00011100101] = 16'b1001110010001110;
	exp_table[11'b00011100110] = 16'b1001110100101011;
	exp_table[11'b00011100111] = 16'b1001110111001000;
	exp_table[11'b00011101000] = 16'b1001111001100110;
	exp_table[11'b00011101001] = 16'b1001111100000101;
	exp_table[11'b00011101010] = 16'b1001111110100100;
	exp_table[11'b00011101011] = 16'b1010000001000100;
	exp_table[11'b00011101100] = 16'b1010000011100101;
	exp_table[11'b00011101101] = 16'b1010000110000110;
	exp_table[11'b00011101110] = 16'b1010001000101000;
	exp_table[11'b00011101111] = 16'b1010001011001010;
	exp_table[11'b00011110000] = 16'b1010001101101110;
	exp_table[11'b00011110001] = 16'b1010010000010001;
	exp_table[11'b00011110010] = 16'b1010010010110110;
	exp_table[11'b00011110011] = 16'b1010010101011011;
	exp_table[11'b00011110100] = 16'b1010011000000000;
	exp_table[11'b00011110101] = 16'b1010011010100111;
	exp_table[11'b00011110110] = 16'b1010011101001110;
	exp_table[11'b00011110111] = 16'b1010011111110101;
	exp_table[11'b00011111000] = 16'b1010100010011110;
	exp_table[11'b00011111001] = 16'b1010100101000111;
	exp_table[11'b00011111010] = 16'b1010100111110000;
	exp_table[11'b00011111011] = 16'b1010101010011010;
	exp_table[11'b00011111100] = 16'b1010101101000101;
	exp_table[11'b00011111101] = 16'b1010101111110001;
	exp_table[11'b00011111110] = 16'b1010110010011101;
	exp_table[11'b00011111111] = 16'b1010110101001010;
	exp_table[11'b00100000000] = 16'b1010110111111000;
	exp_table[11'b00100000001] = 16'b1010111010100110;
	exp_table[11'b00100000010] = 16'b1010111101010101;
	exp_table[11'b00100000011] = 16'b1011000000000101;
	exp_table[11'b00100000100] = 16'b1011000010110101;
	exp_table[11'b00100000101] = 16'b1011000101100110;
	exp_table[11'b00100000110] = 16'b1011001000011000;
	exp_table[11'b00100000111] = 16'b1011001011001010;
	exp_table[11'b00100001000] = 16'b1011001101111110;
	exp_table[11'b00100001001] = 16'b1011010000110001;
	exp_table[11'b00100001010] = 16'b1011010011100110;
	exp_table[11'b00100001011] = 16'b1011010110011011;
	exp_table[11'b00100001100] = 16'b1011011001010001;
	exp_table[11'b00100001101] = 16'b1011011100001000;
	exp_table[11'b00100001110] = 16'b1011011110111111;
	exp_table[11'b00100001111] = 16'b1011100001110111;
	exp_table[11'b00100010000] = 16'b1011100100110000;
	exp_table[11'b00100010001] = 16'b1011100111101010;
	exp_table[11'b00100010010] = 16'b1011101010100100;
	exp_table[11'b00100010011] = 16'b1011101101011111;
	exp_table[11'b00100010100] = 16'b1011110000011011;
	exp_table[11'b00100010101] = 16'b1011110011010111;
	exp_table[11'b00100010110] = 16'b1011110110010100;
	exp_table[11'b00100010111] = 16'b1011111001010010;
	exp_table[11'b00100011000] = 16'b1011111100010001;
	exp_table[11'b00100011001] = 16'b1011111111010001;
	exp_table[11'b00100011010] = 16'b1100000010010001;
	exp_table[11'b00100011011] = 16'b1100000101010010;
	exp_table[11'b00100011100] = 16'b1100001000010011;
	exp_table[11'b00100011101] = 16'b1100001011010110;
	exp_table[11'b00100011110] = 16'b1100001110011001;
	exp_table[11'b00100011111] = 16'b1100010001011101;
	exp_table[11'b00100100000] = 16'b1100010100100010;
	exp_table[11'b00100100001] = 16'b1100010111100111;
	exp_table[11'b00100100010] = 16'b1100011010101110;
	exp_table[11'b00100100011] = 16'b1100011101110101;
	exp_table[11'b00100100100] = 16'b1100100000111101;
	exp_table[11'b00100100101] = 16'b1100100100000101;
	exp_table[11'b00100100110] = 16'b1100100111001111;
	exp_table[11'b00100100111] = 16'b1100101010011001;
	exp_table[11'b00100101000] = 16'b1100101101100100;
	exp_table[11'b00100101001] = 16'b1100110000110000;
	exp_table[11'b00100101010] = 16'b1100110011111100;
	exp_table[11'b00100101011] = 16'b1100110111001010;
	exp_table[11'b00100101100] = 16'b1100111010011000;
	exp_table[11'b00100101101] = 16'b1100111101100111;
	exp_table[11'b00100101110] = 16'b1101000000110111;
	exp_table[11'b00100101111] = 16'b1101000100000111;
	exp_table[11'b00100110000] = 16'b1101000111011001;
	exp_table[11'b00100110001] = 16'b1101001010101011;
	exp_table[11'b00100110010] = 16'b1101001101111110;
	exp_table[11'b00100110011] = 16'b1101010001010010;
	exp_table[11'b00100110100] = 16'b1101010100100111;
	exp_table[11'b00100110101] = 16'b1101010111111100;
	exp_table[11'b00100110110] = 16'b1101011011010011;
	exp_table[11'b00100110111] = 16'b1101011110101010;
	exp_table[11'b00100111000] = 16'b1101100010000010;
	exp_table[11'b00100111001] = 16'b1101100101011011;
	exp_table[11'b00100111010] = 16'b1101101000110101;
	exp_table[11'b00100111011] = 16'b1101101100001111;
	exp_table[11'b00100111100] = 16'b1101101111101011;
	exp_table[11'b00100111101] = 16'b1101110011000111;
	exp_table[11'b00100111110] = 16'b1101110110100100;
	exp_table[11'b00100111111] = 16'b1101111010000010;
	exp_table[11'b00101000000] = 16'b1101111101100001;
	exp_table[11'b00101000001] = 16'b1110000001000001;
	exp_table[11'b00101000010] = 16'b1110000100100010;
	exp_table[11'b00101000011] = 16'b1110001000000011;
	exp_table[11'b00101000100] = 16'b1110001011100110;
	exp_table[11'b00101000101] = 16'b1110001111001001;
	exp_table[11'b00101000110] = 16'b1110010010101101;
	exp_table[11'b00101000111] = 16'b1110010110010011;
	exp_table[11'b00101001000] = 16'b1110011001111001;
	exp_table[11'b00101001001] = 16'b1110011101011111;
	exp_table[11'b00101001010] = 16'b1110100001000111;
	exp_table[11'b00101001011] = 16'b1110100100110000;
	exp_table[11'b00101001100] = 16'b1110101000011010;
	exp_table[11'b00101001101] = 16'b1110101100000100;
	exp_table[11'b00101001110] = 16'b1110101111110000;
	exp_table[11'b00101001111] = 16'b1110110011011100;
	exp_table[11'b00101010000] = 16'b1110110111001001;
	exp_table[11'b00101010001] = 16'b1110111010111000;
	exp_table[11'b00101010010] = 16'b1110111110100111;
	exp_table[11'b00101010011] = 16'b1111000010010111;
	exp_table[11'b00101010100] = 16'b1111000110001000;
	exp_table[11'b00101010101] = 16'b1111001001111010;
	exp_table[11'b00101010110] = 16'b1111001101101101;
	exp_table[11'b00101010111] = 16'b1111010001100001;
	exp_table[11'b00101011000] = 16'b1111010101010110;
	exp_table[11'b00101011001] = 16'b1111011001001100;
	exp_table[11'b00101011010] = 16'b1111011101000010;
	exp_table[11'b00101011011] = 16'b1111100000111010;
	exp_table[11'b00101011100] = 16'b1111100100110011;
	exp_table[11'b00101011101] = 16'b1111101000101101;
	exp_table[11'b00101011110] = 16'b1111101100100111;
	exp_table[11'b00101011111] = 16'b1111110000100011;
	exp_table[11'b00101100000] = 16'b1111110100011111;
	exp_table[11'b00101100001] = 16'b1111111000011101;
	exp_table[11'b00101100010] = 16'b1111111100011100;
	exp_table[11'b00101100011] = 16'b1111111111111111;
	exp_table[11'b00101100100] = 16'b1111111111111111;
	exp_table[11'b00101100101] = 16'b1111111111111111;
	exp_table[11'b00101100110] = 16'b1111111111111111;
	exp_table[11'b00101100111] = 16'b1111111111111111;
	exp_table[11'b00101101000] = 16'b1111111111111111;
	exp_table[11'b00101101001] = 16'b1111111111111111;
	exp_table[11'b00101101010] = 16'b1111111111111111;
	exp_table[11'b00101101011] = 16'b1111111111111111;
	exp_table[11'b00101101100] = 16'b1111111111111111;
	exp_table[11'b00101101101] = 16'b1111111111111111;
	exp_table[11'b00101101110] = 16'b1111111111111111;
	exp_table[11'b00101101111] = 16'b1111111111111111;
	exp_table[11'b00101110000] = 16'b1111111111111111;
	exp_table[11'b00101110001] = 16'b1111111111111111;
	exp_table[11'b00101110010] = 16'b1111111111111111;
	exp_table[11'b00101110011] = 16'b1111111111111111;
	exp_table[11'b00101110100] = 16'b1111111111111111;
	exp_table[11'b00101110101] = 16'b1111111111111111;
	exp_table[11'b00101110110] = 16'b1111111111111111;
	exp_table[11'b00101110111] = 16'b1111111111111111;
	exp_table[11'b00101111000] = 16'b1111111111111111;
	exp_table[11'b00101111001] = 16'b1111111111111111;
	exp_table[11'b00101111010] = 16'b1111111111111111;
	exp_table[11'b00101111011] = 16'b1111111111111111;
	exp_table[11'b00101111100] = 16'b1111111111111111;
	exp_table[11'b00101111101] = 16'b1111111111111111;
	exp_table[11'b00101111110] = 16'b1111111111111111;
	exp_table[11'b00101111111] = 16'b1111111111111111;
	exp_table[11'b00110000000] = 16'b1111111111111111;
	exp_table[11'b00110000001] = 16'b1111111111111111;
	exp_table[11'b00110000010] = 16'b1111111111111111;
	exp_table[11'b00110000011] = 16'b1111111111111111;
	exp_table[11'b00110000100] = 16'b1111111111111111;
	exp_table[11'b00110000101] = 16'b1111111111111111;
	exp_table[11'b00110000110] = 16'b1111111111111111;
	exp_table[11'b00110000111] = 16'b1111111111111111;
	exp_table[11'b00110001000] = 16'b1111111111111111;
	exp_table[11'b00110001001] = 16'b1111111111111111;
	exp_table[11'b00110001010] = 16'b1111111111111111;
	exp_table[11'b00110001011] = 16'b1111111111111111;
	exp_table[11'b00110001100] = 16'b1111111111111111;
	exp_table[11'b00110001101] = 16'b1111111111111111;
	exp_table[11'b00110001110] = 16'b1111111111111111;
	exp_table[11'b00110001111] = 16'b1111111111111111;
	exp_table[11'b00110010000] = 16'b1111111111111111;
	exp_table[11'b00110010001] = 16'b1111111111111111;
	exp_table[11'b00110010010] = 16'b1111111111111111;
	exp_table[11'b00110010011] = 16'b1111111111111111;
	exp_table[11'b00110010100] = 16'b1111111111111111;
	exp_table[11'b00110010101] = 16'b1111111111111111;
	exp_table[11'b00110010110] = 16'b1111111111111111;
	exp_table[11'b00110010111] = 16'b1111111111111111;
	exp_table[11'b00110011000] = 16'b1111111111111111;
	exp_table[11'b00110011001] = 16'b1111111111111111;
	exp_table[11'b00110011010] = 16'b1111111111111111;
	exp_table[11'b00110011011] = 16'b1111111111111111;
	exp_table[11'b00110011100] = 16'b1111111111111111;
	exp_table[11'b00110011101] = 16'b1111111111111111;
	exp_table[11'b00110011110] = 16'b1111111111111111;
	exp_table[11'b00110011111] = 16'b1111111111111111;
	exp_table[11'b00110100000] = 16'b1111111111111111;
	exp_table[11'b00110100001] = 16'b1111111111111111;
	exp_table[11'b00110100010] = 16'b1111111111111111;
	exp_table[11'b00110100011] = 16'b1111111111111111;
	exp_table[11'b00110100100] = 16'b1111111111111111;
	exp_table[11'b00110100101] = 16'b1111111111111111;
	exp_table[11'b00110100110] = 16'b1111111111111111;
	exp_table[11'b00110100111] = 16'b1111111111111111;
	exp_table[11'b00110101000] = 16'b1111111111111111;
	exp_table[11'b00110101001] = 16'b1111111111111111;
	exp_table[11'b00110101010] = 16'b1111111111111111;
	exp_table[11'b00110101011] = 16'b1111111111111111;
	exp_table[11'b00110101100] = 16'b1111111111111111;
	exp_table[11'b00110101101] = 16'b1111111111111111;
	exp_table[11'b00110101110] = 16'b1111111111111111;
	exp_table[11'b00110101111] = 16'b1111111111111111;
	exp_table[11'b00110110000] = 16'b1111111111111111;
	exp_table[11'b00110110001] = 16'b1111111111111111;
	exp_table[11'b00110110010] = 16'b1111111111111111;
	exp_table[11'b00110110011] = 16'b1111111111111111;
	exp_table[11'b00110110100] = 16'b1111111111111111;
	exp_table[11'b00110110101] = 16'b1111111111111111;
	exp_table[11'b00110110110] = 16'b1111111111111111;
	exp_table[11'b00110110111] = 16'b1111111111111111;
	exp_table[11'b00110111000] = 16'b1111111111111111;
	exp_table[11'b00110111001] = 16'b1111111111111111;
	exp_table[11'b00110111010] = 16'b1111111111111111;
	exp_table[11'b00110111011] = 16'b1111111111111111;
	exp_table[11'b00110111100] = 16'b1111111111111111;
	exp_table[11'b00110111101] = 16'b1111111111111111;
	exp_table[11'b00110111110] = 16'b1111111111111111;
	exp_table[11'b00110111111] = 16'b1111111111111111;
	exp_table[11'b00111000000] = 16'b1111111111111111;
	exp_table[11'b00111000001] = 16'b1111111111111111;
	exp_table[11'b00111000010] = 16'b1111111111111111;
	exp_table[11'b00111000011] = 16'b1111111111111111;
	exp_table[11'b00111000100] = 16'b1111111111111111;
	exp_table[11'b00111000101] = 16'b1111111111111111;
	exp_table[11'b00111000110] = 16'b1111111111111111;
	exp_table[11'b00111000111] = 16'b1111111111111111;
	exp_table[11'b00111001000] = 16'b1111111111111111;
	exp_table[11'b00111001001] = 16'b1111111111111111;
	exp_table[11'b00111001010] = 16'b1111111111111111;
	exp_table[11'b00111001011] = 16'b1111111111111111;
	exp_table[11'b00111001100] = 16'b1111111111111111;
	exp_table[11'b00111001101] = 16'b1111111111111111;
	exp_table[11'b00111001110] = 16'b1111111111111111;
	exp_table[11'b00111001111] = 16'b1111111111111111;
	exp_table[11'b00111010000] = 16'b1111111111111111;
	exp_table[11'b00111010001] = 16'b1111111111111111;
	exp_table[11'b00111010010] = 16'b1111111111111111;
	exp_table[11'b00111010011] = 16'b1111111111111111;
	exp_table[11'b00111010100] = 16'b1111111111111111;
	exp_table[11'b00111010101] = 16'b1111111111111111;
	exp_table[11'b00111010110] = 16'b1111111111111111;
	exp_table[11'b00111010111] = 16'b1111111111111111;
	exp_table[11'b00111011000] = 16'b1111111111111111;
	exp_table[11'b00111011001] = 16'b1111111111111111;
	exp_table[11'b00111011010] = 16'b1111111111111111;
	exp_table[11'b00111011011] = 16'b1111111111111111;
	exp_table[11'b00111011100] = 16'b1111111111111111;
	exp_table[11'b00111011101] = 16'b1111111111111111;
	exp_table[11'b00111011110] = 16'b1111111111111111;
	exp_table[11'b00111011111] = 16'b1111111111111111;
	exp_table[11'b00111100000] = 16'b1111111111111111;
	exp_table[11'b00111100001] = 16'b1111111111111111;
	exp_table[11'b00111100010] = 16'b1111111111111111;
	exp_table[11'b00111100011] = 16'b1111111111111111;
	exp_table[11'b00111100100] = 16'b1111111111111111;
	exp_table[11'b00111100101] = 16'b1111111111111111;
	exp_table[11'b00111100110] = 16'b1111111111111111;
	exp_table[11'b00111100111] = 16'b1111111111111111;
	exp_table[11'b00111101000] = 16'b1111111111111111;
	exp_table[11'b00111101001] = 16'b1111111111111111;
	exp_table[11'b00111101010] = 16'b1111111111111111;
	exp_table[11'b00111101011] = 16'b1111111111111111;
	exp_table[11'b00111101100] = 16'b1111111111111111;
	exp_table[11'b00111101101] = 16'b1111111111111111;
	exp_table[11'b00111101110] = 16'b1111111111111111;
	exp_table[11'b00111101111] = 16'b1111111111111111;
	exp_table[11'b00111110000] = 16'b1111111111111111;
	exp_table[11'b00111110001] = 16'b1111111111111111;
	exp_table[11'b00111110010] = 16'b1111111111111111;
	exp_table[11'b00111110011] = 16'b1111111111111111;
	exp_table[11'b00111110100] = 16'b1111111111111111;
	exp_table[11'b00111110101] = 16'b1111111111111111;
	exp_table[11'b00111110110] = 16'b1111111111111111;
	exp_table[11'b00111110111] = 16'b1111111111111111;
	exp_table[11'b00111111000] = 16'b1111111111111111;
	exp_table[11'b00111111001] = 16'b1111111111111111;
	exp_table[11'b00111111010] = 16'b1111111111111111;
	exp_table[11'b00111111011] = 16'b1111111111111111;
	exp_table[11'b00111111100] = 16'b1111111111111111;
	exp_table[11'b00111111101] = 16'b1111111111111111;
	exp_table[11'b00111111110] = 16'b1111111111111111;
	exp_table[11'b00111111111] = 16'b1111111111111111;
	exp_table[11'b01000000000] = 16'b1111111111111111;
	exp_table[11'b01000000001] = 16'b1111111111111111;
	exp_table[11'b01000000010] = 16'b1111111111111111;
	exp_table[11'b01000000011] = 16'b1111111111111111;
	exp_table[11'b01000000100] = 16'b1111111111111111;
	exp_table[11'b01000000101] = 16'b1111111111111111;
	exp_table[11'b01000000110] = 16'b1111111111111111;
	exp_table[11'b01000000111] = 16'b1111111111111111;
	exp_table[11'b01000001000] = 16'b1111111111111111;
	exp_table[11'b01000001001] = 16'b1111111111111111;
	exp_table[11'b01000001010] = 16'b1111111111111111;
	exp_table[11'b01000001011] = 16'b1111111111111111;
	exp_table[11'b01000001100] = 16'b1111111111111111;
	exp_table[11'b01000001101] = 16'b1111111111111111;
	exp_table[11'b01000001110] = 16'b1111111111111111;
	exp_table[11'b01000001111] = 16'b1111111111111111;
	exp_table[11'b01000010000] = 16'b1111111111111111;
	exp_table[11'b01000010001] = 16'b1111111111111111;
	exp_table[11'b01000010010] = 16'b1111111111111111;
	exp_table[11'b01000010011] = 16'b1111111111111111;
	exp_table[11'b01000010100] = 16'b1111111111111111;
	exp_table[11'b01000010101] = 16'b1111111111111111;
	exp_table[11'b01000010110] = 16'b1111111111111111;
	exp_table[11'b01000010111] = 16'b1111111111111111;
	exp_table[11'b01000011000] = 16'b1111111111111111;
	exp_table[11'b01000011001] = 16'b1111111111111111;
	exp_table[11'b01000011010] = 16'b1111111111111111;
	exp_table[11'b01000011011] = 16'b1111111111111111;
	exp_table[11'b01000011100] = 16'b1111111111111111;
	exp_table[11'b01000011101] = 16'b1111111111111111;
	exp_table[11'b01000011110] = 16'b1111111111111111;
	exp_table[11'b01000011111] = 16'b1111111111111111;
	exp_table[11'b01000100000] = 16'b1111111111111111;
	exp_table[11'b01000100001] = 16'b1111111111111111;
	exp_table[11'b01000100010] = 16'b1111111111111111;
	exp_table[11'b01000100011] = 16'b1111111111111111;
	exp_table[11'b01000100100] = 16'b1111111111111111;
	exp_table[11'b01000100101] = 16'b1111111111111111;
	exp_table[11'b01000100110] = 16'b1111111111111111;
	exp_table[11'b01000100111] = 16'b1111111111111111;
	exp_table[11'b01000101000] = 16'b1111111111111111;
	exp_table[11'b01000101001] = 16'b1111111111111111;
	exp_table[11'b01000101010] = 16'b1111111111111111;
	exp_table[11'b01000101011] = 16'b1111111111111111;
	exp_table[11'b01000101100] = 16'b1111111111111111;
	exp_table[11'b01000101101] = 16'b1111111111111111;
	exp_table[11'b01000101110] = 16'b1111111111111111;
	exp_table[11'b01000101111] = 16'b1111111111111111;
	exp_table[11'b01000110000] = 16'b1111111111111111;
	exp_table[11'b01000110001] = 16'b1111111111111111;
	exp_table[11'b01000110010] = 16'b1111111111111111;
	exp_table[11'b01000110011] = 16'b1111111111111111;
	exp_table[11'b01000110100] = 16'b1111111111111111;
	exp_table[11'b01000110101] = 16'b1111111111111111;
	exp_table[11'b01000110110] = 16'b1111111111111111;
	exp_table[11'b01000110111] = 16'b1111111111111111;
	exp_table[11'b01000111000] = 16'b1111111111111111;
	exp_table[11'b01000111001] = 16'b1111111111111111;
	exp_table[11'b01000111010] = 16'b1111111111111111;
	exp_table[11'b01000111011] = 16'b1111111111111111;
	exp_table[11'b01000111100] = 16'b1111111111111111;
	exp_table[11'b01000111101] = 16'b1111111111111111;
	exp_table[11'b01000111110] = 16'b1111111111111111;
	exp_table[11'b01000111111] = 16'b1111111111111111;
	exp_table[11'b01001000000] = 16'b1111111111111111;
	exp_table[11'b01001000001] = 16'b1111111111111111;
	exp_table[11'b01001000010] = 16'b1111111111111111;
	exp_table[11'b01001000011] = 16'b1111111111111111;
	exp_table[11'b01001000100] = 16'b1111111111111111;
	exp_table[11'b01001000101] = 16'b1111111111111111;
	exp_table[11'b01001000110] = 16'b1111111111111111;
	exp_table[11'b01001000111] = 16'b1111111111111111;
	exp_table[11'b01001001000] = 16'b1111111111111111;
	exp_table[11'b01001001001] = 16'b1111111111111111;
	exp_table[11'b01001001010] = 16'b1111111111111111;
	exp_table[11'b01001001011] = 16'b1111111111111111;
	exp_table[11'b01001001100] = 16'b1111111111111111;
	exp_table[11'b01001001101] = 16'b1111111111111111;
	exp_table[11'b01001001110] = 16'b1111111111111111;
	exp_table[11'b01001001111] = 16'b1111111111111111;
	exp_table[11'b01001010000] = 16'b1111111111111111;
	exp_table[11'b01001010001] = 16'b1111111111111111;
	exp_table[11'b01001010010] = 16'b1111111111111111;
	exp_table[11'b01001010011] = 16'b1111111111111111;
	exp_table[11'b01001010100] = 16'b1111111111111111;
	exp_table[11'b01001010101] = 16'b1111111111111111;
	exp_table[11'b01001010110] = 16'b1111111111111111;
	exp_table[11'b01001010111] = 16'b1111111111111111;
	exp_table[11'b01001011000] = 16'b1111111111111111;
	exp_table[11'b01001011001] = 16'b1111111111111111;
	exp_table[11'b01001011010] = 16'b1111111111111111;
	exp_table[11'b01001011011] = 16'b1111111111111111;
	exp_table[11'b01001011100] = 16'b1111111111111111;
	exp_table[11'b01001011101] = 16'b1111111111111111;
	exp_table[11'b01001011110] = 16'b1111111111111111;
	exp_table[11'b01001011111] = 16'b1111111111111111;
	exp_table[11'b01001100000] = 16'b1111111111111111;
	exp_table[11'b01001100001] = 16'b1111111111111111;
	exp_table[11'b01001100010] = 16'b1111111111111111;
	exp_table[11'b01001100011] = 16'b1111111111111111;
	exp_table[11'b01001100100] = 16'b1111111111111111;
	exp_table[11'b01001100101] = 16'b1111111111111111;
	exp_table[11'b01001100110] = 16'b1111111111111111;
	exp_table[11'b01001100111] = 16'b1111111111111111;
	exp_table[11'b01001101000] = 16'b1111111111111111;
	exp_table[11'b01001101001] = 16'b1111111111111111;
	exp_table[11'b01001101010] = 16'b1111111111111111;
	exp_table[11'b01001101011] = 16'b1111111111111111;
	exp_table[11'b01001101100] = 16'b1111111111111111;
	exp_table[11'b01001101101] = 16'b1111111111111111;
	exp_table[11'b01001101110] = 16'b1111111111111111;
	exp_table[11'b01001101111] = 16'b1111111111111111;
	exp_table[11'b01001110000] = 16'b1111111111111111;
	exp_table[11'b01001110001] = 16'b1111111111111111;
	exp_table[11'b01001110010] = 16'b1111111111111111;
	exp_table[11'b01001110011] = 16'b1111111111111111;
	exp_table[11'b01001110100] = 16'b1111111111111111;
	exp_table[11'b01001110101] = 16'b1111111111111111;
	exp_table[11'b01001110110] = 16'b1111111111111111;
	exp_table[11'b01001110111] = 16'b1111111111111111;
	exp_table[11'b01001111000] = 16'b1111111111111111;
	exp_table[11'b01001111001] = 16'b1111111111111111;
	exp_table[11'b01001111010] = 16'b1111111111111111;
	exp_table[11'b01001111011] = 16'b1111111111111111;
	exp_table[11'b01001111100] = 16'b1111111111111111;
	exp_table[11'b01001111101] = 16'b1111111111111111;
	exp_table[11'b01001111110] = 16'b1111111111111111;
	exp_table[11'b01001111111] = 16'b1111111111111111;
	exp_table[11'b01010000000] = 16'b1111111111111111;
	exp_table[11'b01010000001] = 16'b1111111111111111;
	exp_table[11'b01010000010] = 16'b1111111111111111;
	exp_table[11'b01010000011] = 16'b1111111111111111;
	exp_table[11'b01010000100] = 16'b1111111111111111;
	exp_table[11'b01010000101] = 16'b1111111111111111;
	exp_table[11'b01010000110] = 16'b1111111111111111;
	exp_table[11'b01010000111] = 16'b1111111111111111;
	exp_table[11'b01010001000] = 16'b1111111111111111;
	exp_table[11'b01010001001] = 16'b1111111111111111;
	exp_table[11'b01010001010] = 16'b1111111111111111;
	exp_table[11'b01010001011] = 16'b1111111111111111;
	exp_table[11'b01010001100] = 16'b1111111111111111;
	exp_table[11'b01010001101] = 16'b1111111111111111;
	exp_table[11'b01010001110] = 16'b1111111111111111;
	exp_table[11'b01010001111] = 16'b1111111111111111;
	exp_table[11'b01010010000] = 16'b1111111111111111;
	exp_table[11'b01010010001] = 16'b1111111111111111;
	exp_table[11'b01010010010] = 16'b1111111111111111;
	exp_table[11'b01010010011] = 16'b1111111111111111;
	exp_table[11'b01010010100] = 16'b1111111111111111;
	exp_table[11'b01010010101] = 16'b1111111111111111;
	exp_table[11'b01010010110] = 16'b1111111111111111;
	exp_table[11'b01010010111] = 16'b1111111111111111;
	exp_table[11'b01010011000] = 16'b1111111111111111;
	exp_table[11'b01010011001] = 16'b1111111111111111;
	exp_table[11'b01010011010] = 16'b1111111111111111;
	exp_table[11'b01010011011] = 16'b1111111111111111;
	exp_table[11'b01010011100] = 16'b1111111111111111;
	exp_table[11'b01010011101] = 16'b1111111111111111;
	exp_table[11'b01010011110] = 16'b1111111111111111;
	exp_table[11'b01010011111] = 16'b1111111111111111;
	exp_table[11'b01010100000] = 16'b1111111111111111;
	exp_table[11'b01010100001] = 16'b1111111111111111;
	exp_table[11'b01010100010] = 16'b1111111111111111;
	exp_table[11'b01010100011] = 16'b1111111111111111;
	exp_table[11'b01010100100] = 16'b1111111111111111;
	exp_table[11'b01010100101] = 16'b1111111111111111;
	exp_table[11'b01010100110] = 16'b1111111111111111;
	exp_table[11'b01010100111] = 16'b1111111111111111;
	exp_table[11'b01010101000] = 16'b1111111111111111;
	exp_table[11'b01010101001] = 16'b1111111111111111;
	exp_table[11'b01010101010] = 16'b1111111111111111;
	exp_table[11'b01010101011] = 16'b1111111111111111;
	exp_table[11'b01010101100] = 16'b1111111111111111;
	exp_table[11'b01010101101] = 16'b1111111111111111;
	exp_table[11'b01010101110] = 16'b1111111111111111;
	exp_table[11'b01010101111] = 16'b1111111111111111;
	exp_table[11'b01010110000] = 16'b1111111111111111;
	exp_table[11'b01010110001] = 16'b1111111111111111;
	exp_table[11'b01010110010] = 16'b1111111111111111;
	exp_table[11'b01010110011] = 16'b1111111111111111;
	exp_table[11'b01010110100] = 16'b1111111111111111;
	exp_table[11'b01010110101] = 16'b1111111111111111;
	exp_table[11'b01010110110] = 16'b1111111111111111;
	exp_table[11'b01010110111] = 16'b1111111111111111;
	exp_table[11'b01010111000] = 16'b1111111111111111;
	exp_table[11'b01010111001] = 16'b1111111111111111;
	exp_table[11'b01010111010] = 16'b1111111111111111;
	exp_table[11'b01010111011] = 16'b1111111111111111;
	exp_table[11'b01010111100] = 16'b1111111111111111;
	exp_table[11'b01010111101] = 16'b1111111111111111;
	exp_table[11'b01010111110] = 16'b1111111111111111;
	exp_table[11'b01010111111] = 16'b1111111111111111;
	exp_table[11'b01011000000] = 16'b1111111111111111;
	exp_table[11'b01011000001] = 16'b1111111111111111;
	exp_table[11'b01011000010] = 16'b1111111111111111;
	exp_table[11'b01011000011] = 16'b1111111111111111;
	exp_table[11'b01011000100] = 16'b1111111111111111;
	exp_table[11'b01011000101] = 16'b1111111111111111;
	exp_table[11'b01011000110] = 16'b1111111111111111;
	exp_table[11'b01011000111] = 16'b1111111111111111;
	exp_table[11'b01011001000] = 16'b1111111111111111;
	exp_table[11'b01011001001] = 16'b1111111111111111;
	exp_table[11'b01011001010] = 16'b1111111111111111;
	exp_table[11'b01011001011] = 16'b1111111111111111;
	exp_table[11'b01011001100] = 16'b1111111111111111;
	exp_table[11'b01011001101] = 16'b1111111111111111;
	exp_table[11'b01011001110] = 16'b1111111111111111;
	exp_table[11'b01011001111] = 16'b1111111111111111;
	exp_table[11'b01011010000] = 16'b1111111111111111;
	exp_table[11'b01011010001] = 16'b1111111111111111;
	exp_table[11'b01011010010] = 16'b1111111111111111;
	exp_table[11'b01011010011] = 16'b1111111111111111;
	exp_table[11'b01011010100] = 16'b1111111111111111;
	exp_table[11'b01011010101] = 16'b1111111111111111;
	exp_table[11'b01011010110] = 16'b1111111111111111;
	exp_table[11'b01011010111] = 16'b1111111111111111;
	exp_table[11'b01011011000] = 16'b1111111111111111;
	exp_table[11'b01011011001] = 16'b1111111111111111;
	exp_table[11'b01011011010] = 16'b1111111111111111;
	exp_table[11'b01011011011] = 16'b1111111111111111;
	exp_table[11'b01011011100] = 16'b1111111111111111;
	exp_table[11'b01011011101] = 16'b1111111111111111;
	exp_table[11'b01011011110] = 16'b1111111111111111;
	exp_table[11'b01011011111] = 16'b1111111111111111;
	exp_table[11'b01011100000] = 16'b1111111111111111;
	exp_table[11'b01011100001] = 16'b1111111111111111;
	exp_table[11'b01011100010] = 16'b1111111111111111;
	exp_table[11'b01011100011] = 16'b1111111111111111;
	exp_table[11'b01011100100] = 16'b1111111111111111;
	exp_table[11'b01011100101] = 16'b1111111111111111;
	exp_table[11'b01011100110] = 16'b1111111111111111;
	exp_table[11'b01011100111] = 16'b1111111111111111;
	exp_table[11'b01011101000] = 16'b1111111111111111;
	exp_table[11'b01011101001] = 16'b1111111111111111;
	exp_table[11'b01011101010] = 16'b1111111111111111;
	exp_table[11'b01011101011] = 16'b1111111111111111;
	exp_table[11'b01011101100] = 16'b1111111111111111;
	exp_table[11'b01011101101] = 16'b1111111111111111;
	exp_table[11'b01011101110] = 16'b1111111111111111;
	exp_table[11'b01011101111] = 16'b1111111111111111;
	exp_table[11'b01011110000] = 16'b1111111111111111;
	exp_table[11'b01011110001] = 16'b1111111111111111;
	exp_table[11'b01011110010] = 16'b1111111111111111;
	exp_table[11'b01011110011] = 16'b1111111111111111;
	exp_table[11'b01011110100] = 16'b1111111111111111;
	exp_table[11'b01011110101] = 16'b1111111111111111;
	exp_table[11'b01011110110] = 16'b1111111111111111;
	exp_table[11'b01011110111] = 16'b1111111111111111;
	exp_table[11'b01011111000] = 16'b1111111111111111;
	exp_table[11'b01011111001] = 16'b1111111111111111;
	exp_table[11'b01011111010] = 16'b1111111111111111;
	exp_table[11'b01011111011] = 16'b1111111111111111;
	exp_table[11'b01011111100] = 16'b1111111111111111;
	exp_table[11'b01011111101] = 16'b1111111111111111;
	exp_table[11'b01011111110] = 16'b1111111111111111;
	exp_table[11'b01011111111] = 16'b1111111111111111;
	exp_table[11'b01100000000] = 16'b1111111111111111;
	exp_table[11'b01100000001] = 16'b1111111111111111;
	exp_table[11'b01100000010] = 16'b1111111111111111;
	exp_table[11'b01100000011] = 16'b1111111111111111;
	exp_table[11'b01100000100] = 16'b1111111111111111;
	exp_table[11'b01100000101] = 16'b1111111111111111;
	exp_table[11'b01100000110] = 16'b1111111111111111;
	exp_table[11'b01100000111] = 16'b1111111111111111;
	exp_table[11'b01100001000] = 16'b1111111111111111;
	exp_table[11'b01100001001] = 16'b1111111111111111;
	exp_table[11'b01100001010] = 16'b1111111111111111;
	exp_table[11'b01100001011] = 16'b1111111111111111;
	exp_table[11'b01100001100] = 16'b1111111111111111;
	exp_table[11'b01100001101] = 16'b1111111111111111;
	exp_table[11'b01100001110] = 16'b1111111111111111;
	exp_table[11'b01100001111] = 16'b1111111111111111;
	exp_table[11'b01100010000] = 16'b1111111111111111;
	exp_table[11'b01100010001] = 16'b1111111111111111;
	exp_table[11'b01100010010] = 16'b1111111111111111;
	exp_table[11'b01100010011] = 16'b1111111111111111;
	exp_table[11'b01100010100] = 16'b1111111111111111;
	exp_table[11'b01100010101] = 16'b1111111111111111;
	exp_table[11'b01100010110] = 16'b1111111111111111;
	exp_table[11'b01100010111] = 16'b1111111111111111;
	exp_table[11'b01100011000] = 16'b1111111111111111;
	exp_table[11'b01100011001] = 16'b1111111111111111;
	exp_table[11'b01100011010] = 16'b1111111111111111;
	exp_table[11'b01100011011] = 16'b1111111111111111;
	exp_table[11'b01100011100] = 16'b1111111111111111;
	exp_table[11'b01100011101] = 16'b1111111111111111;
	exp_table[11'b01100011110] = 16'b1111111111111111;
	exp_table[11'b01100011111] = 16'b1111111111111111;
	exp_table[11'b01100100000] = 16'b1111111111111111;
	exp_table[11'b01100100001] = 16'b1111111111111111;
	exp_table[11'b01100100010] = 16'b1111111111111111;
	exp_table[11'b01100100011] = 16'b1111111111111111;
	exp_table[11'b01100100100] = 16'b1111111111111111;
	exp_table[11'b01100100101] = 16'b1111111111111111;
	exp_table[11'b01100100110] = 16'b1111111111111111;
	exp_table[11'b01100100111] = 16'b1111111111111111;
	exp_table[11'b01100101000] = 16'b1111111111111111;
	exp_table[11'b01100101001] = 16'b1111111111111111;
	exp_table[11'b01100101010] = 16'b1111111111111111;
	exp_table[11'b01100101011] = 16'b1111111111111111;
	exp_table[11'b01100101100] = 16'b1111111111111111;
	exp_table[11'b01100101101] = 16'b1111111111111111;
	exp_table[11'b01100101110] = 16'b1111111111111111;
	exp_table[11'b01100101111] = 16'b1111111111111111;
	exp_table[11'b01100110000] = 16'b1111111111111111;
	exp_table[11'b01100110001] = 16'b1111111111111111;
	exp_table[11'b01100110010] = 16'b1111111111111111;
	exp_table[11'b01100110011] = 16'b1111111111111111;
	exp_table[11'b01100110100] = 16'b1111111111111111;
	exp_table[11'b01100110101] = 16'b1111111111111111;
	exp_table[11'b01100110110] = 16'b1111111111111111;
	exp_table[11'b01100110111] = 16'b1111111111111111;
	exp_table[11'b01100111000] = 16'b1111111111111111;
	exp_table[11'b01100111001] = 16'b1111111111111111;
	exp_table[11'b01100111010] = 16'b1111111111111111;
	exp_table[11'b01100111011] = 16'b1111111111111111;
	exp_table[11'b01100111100] = 16'b1111111111111111;
	exp_table[11'b01100111101] = 16'b1111111111111111;
	exp_table[11'b01100111110] = 16'b1111111111111111;
	exp_table[11'b01100111111] = 16'b1111111111111111;
	exp_table[11'b01101000000] = 16'b1111111111111111;
	exp_table[11'b01101000001] = 16'b1111111111111111;
	exp_table[11'b01101000010] = 16'b1111111111111111;
	exp_table[11'b01101000011] = 16'b1111111111111111;
	exp_table[11'b01101000100] = 16'b1111111111111111;
	exp_table[11'b01101000101] = 16'b1111111111111111;
	exp_table[11'b01101000110] = 16'b1111111111111111;
	exp_table[11'b01101000111] = 16'b1111111111111111;
	exp_table[11'b01101001000] = 16'b1111111111111111;
	exp_table[11'b01101001001] = 16'b1111111111111111;
	exp_table[11'b01101001010] = 16'b1111111111111111;
	exp_table[11'b01101001011] = 16'b1111111111111111;
	exp_table[11'b01101001100] = 16'b1111111111111111;
	exp_table[11'b01101001101] = 16'b1111111111111111;
	exp_table[11'b01101001110] = 16'b1111111111111111;
	exp_table[11'b01101001111] = 16'b1111111111111111;
	exp_table[11'b01101010000] = 16'b1111111111111111;
	exp_table[11'b01101010001] = 16'b1111111111111111;
	exp_table[11'b01101010010] = 16'b1111111111111111;
	exp_table[11'b01101010011] = 16'b1111111111111111;
	exp_table[11'b01101010100] = 16'b1111111111111111;
	exp_table[11'b01101010101] = 16'b1111111111111111;
	exp_table[11'b01101010110] = 16'b1111111111111111;
	exp_table[11'b01101010111] = 16'b1111111111111111;
	exp_table[11'b01101011000] = 16'b1111111111111111;
	exp_table[11'b01101011001] = 16'b1111111111111111;
	exp_table[11'b01101011010] = 16'b1111111111111111;
	exp_table[11'b01101011011] = 16'b1111111111111111;
	exp_table[11'b01101011100] = 16'b1111111111111111;
	exp_table[11'b01101011101] = 16'b1111111111111111;
	exp_table[11'b01101011110] = 16'b1111111111111111;
	exp_table[11'b01101011111] = 16'b1111111111111111;
	exp_table[11'b01101100000] = 16'b1111111111111111;
	exp_table[11'b01101100001] = 16'b1111111111111111;
	exp_table[11'b01101100010] = 16'b1111111111111111;
	exp_table[11'b01101100011] = 16'b1111111111111111;
	exp_table[11'b01101100100] = 16'b1111111111111111;
	exp_table[11'b01101100101] = 16'b1111111111111111;
	exp_table[11'b01101100110] = 16'b1111111111111111;
	exp_table[11'b01101100111] = 16'b1111111111111111;
	exp_table[11'b01101101000] = 16'b1111111111111111;
	exp_table[11'b01101101001] = 16'b1111111111111111;
	exp_table[11'b01101101010] = 16'b1111111111111111;
	exp_table[11'b01101101011] = 16'b1111111111111111;
	exp_table[11'b01101101100] = 16'b1111111111111111;
	exp_table[11'b01101101101] = 16'b1111111111111111;
	exp_table[11'b01101101110] = 16'b1111111111111111;
	exp_table[11'b01101101111] = 16'b1111111111111111;
	exp_table[11'b01101110000] = 16'b1111111111111111;
	exp_table[11'b01101110001] = 16'b1111111111111111;
	exp_table[11'b01101110010] = 16'b1111111111111111;
	exp_table[11'b01101110011] = 16'b1111111111111111;
	exp_table[11'b01101110100] = 16'b1111111111111111;
	exp_table[11'b01101110101] = 16'b1111111111111111;
	exp_table[11'b01101110110] = 16'b1111111111111111;
	exp_table[11'b01101110111] = 16'b1111111111111111;
	exp_table[11'b01101111000] = 16'b1111111111111111;
	exp_table[11'b01101111001] = 16'b1111111111111111;
	exp_table[11'b01101111010] = 16'b1111111111111111;
	exp_table[11'b01101111011] = 16'b1111111111111111;
	exp_table[11'b01101111100] = 16'b1111111111111111;
	exp_table[11'b01101111101] = 16'b1111111111111111;
	exp_table[11'b01101111110] = 16'b1111111111111111;
	exp_table[11'b01101111111] = 16'b1111111111111111;
	exp_table[11'b01110000000] = 16'b1111111111111111;
	exp_table[11'b01110000001] = 16'b1111111111111111;
	exp_table[11'b01110000010] = 16'b1111111111111111;
	exp_table[11'b01110000011] = 16'b1111111111111111;
	exp_table[11'b01110000100] = 16'b1111111111111111;
	exp_table[11'b01110000101] = 16'b1111111111111111;
	exp_table[11'b01110000110] = 16'b1111111111111111;
	exp_table[11'b01110000111] = 16'b1111111111111111;
	exp_table[11'b01110001000] = 16'b1111111111111111;
	exp_table[11'b01110001001] = 16'b1111111111111111;
	exp_table[11'b01110001010] = 16'b1111111111111111;
	exp_table[11'b01110001011] = 16'b1111111111111111;
	exp_table[11'b01110001100] = 16'b1111111111111111;
	exp_table[11'b01110001101] = 16'b1111111111111111;
	exp_table[11'b01110001110] = 16'b1111111111111111;
	exp_table[11'b01110001111] = 16'b1111111111111111;
	exp_table[11'b01110010000] = 16'b1111111111111111;
	exp_table[11'b01110010001] = 16'b1111111111111111;
	exp_table[11'b01110010010] = 16'b1111111111111111;
	exp_table[11'b01110010011] = 16'b1111111111111111;
	exp_table[11'b01110010100] = 16'b1111111111111111;
	exp_table[11'b01110010101] = 16'b1111111111111111;
	exp_table[11'b01110010110] = 16'b1111111111111111;
	exp_table[11'b01110010111] = 16'b1111111111111111;
	exp_table[11'b01110011000] = 16'b1111111111111111;
	exp_table[11'b01110011001] = 16'b1111111111111111;
	exp_table[11'b01110011010] = 16'b1111111111111111;
	exp_table[11'b01110011011] = 16'b1111111111111111;
	exp_table[11'b01110011100] = 16'b1111111111111111;
	exp_table[11'b01110011101] = 16'b1111111111111111;
	exp_table[11'b01110011110] = 16'b1111111111111111;
	exp_table[11'b01110011111] = 16'b1111111111111111;
	exp_table[11'b01110100000] = 16'b1111111111111111;
	exp_table[11'b01110100001] = 16'b1111111111111111;
	exp_table[11'b01110100010] = 16'b1111111111111111;
	exp_table[11'b01110100011] = 16'b1111111111111111;
	exp_table[11'b01110100100] = 16'b1111111111111111;
	exp_table[11'b01110100101] = 16'b1111111111111111;
	exp_table[11'b01110100110] = 16'b1111111111111111;
	exp_table[11'b01110100111] = 16'b1111111111111111;
	exp_table[11'b01110101000] = 16'b1111111111111111;
	exp_table[11'b01110101001] = 16'b1111111111111111;
	exp_table[11'b01110101010] = 16'b1111111111111111;
	exp_table[11'b01110101011] = 16'b1111111111111111;
	exp_table[11'b01110101100] = 16'b1111111111111111;
	exp_table[11'b01110101101] = 16'b1111111111111111;
	exp_table[11'b01110101110] = 16'b1111111111111111;
	exp_table[11'b01110101111] = 16'b1111111111111111;
	exp_table[11'b01110110000] = 16'b1111111111111111;
	exp_table[11'b01110110001] = 16'b1111111111111111;
	exp_table[11'b01110110010] = 16'b1111111111111111;
	exp_table[11'b01110110011] = 16'b1111111111111111;
	exp_table[11'b01110110100] = 16'b1111111111111111;
	exp_table[11'b01110110101] = 16'b1111111111111111;
	exp_table[11'b01110110110] = 16'b1111111111111111;
	exp_table[11'b01110110111] = 16'b1111111111111111;
	exp_table[11'b01110111000] = 16'b1111111111111111;
	exp_table[11'b01110111001] = 16'b1111111111111111;
	exp_table[11'b01110111010] = 16'b1111111111111111;
	exp_table[11'b01110111011] = 16'b1111111111111111;
	exp_table[11'b01110111100] = 16'b1111111111111111;
	exp_table[11'b01110111101] = 16'b1111111111111111;
	exp_table[11'b01110111110] = 16'b1111111111111111;
	exp_table[11'b01110111111] = 16'b1111111111111111;
	exp_table[11'b01111000000] = 16'b1111111111111111;
	exp_table[11'b01111000001] = 16'b1111111111111111;
	exp_table[11'b01111000010] = 16'b1111111111111111;
	exp_table[11'b01111000011] = 16'b1111111111111111;
	exp_table[11'b01111000100] = 16'b1111111111111111;
	exp_table[11'b01111000101] = 16'b1111111111111111;
	exp_table[11'b01111000110] = 16'b1111111111111111;
	exp_table[11'b01111000111] = 16'b1111111111111111;
	exp_table[11'b01111001000] = 16'b1111111111111111;
	exp_table[11'b01111001001] = 16'b1111111111111111;
	exp_table[11'b01111001010] = 16'b1111111111111111;
	exp_table[11'b01111001011] = 16'b1111111111111111;
	exp_table[11'b01111001100] = 16'b1111111111111111;
	exp_table[11'b01111001101] = 16'b1111111111111111;
	exp_table[11'b01111001110] = 16'b1111111111111111;
	exp_table[11'b01111001111] = 16'b1111111111111111;
	exp_table[11'b01111010000] = 16'b1111111111111111;
	exp_table[11'b01111010001] = 16'b1111111111111111;
	exp_table[11'b01111010010] = 16'b1111111111111111;
	exp_table[11'b01111010011] = 16'b1111111111111111;
	exp_table[11'b01111010100] = 16'b1111111111111111;
	exp_table[11'b01111010101] = 16'b1111111111111111;
	exp_table[11'b01111010110] = 16'b1111111111111111;
	exp_table[11'b01111010111] = 16'b1111111111111111;
	exp_table[11'b01111011000] = 16'b1111111111111111;
	exp_table[11'b01111011001] = 16'b1111111111111111;
	exp_table[11'b01111011010] = 16'b1111111111111111;
	exp_table[11'b01111011011] = 16'b1111111111111111;
	exp_table[11'b01111011100] = 16'b1111111111111111;
	exp_table[11'b01111011101] = 16'b1111111111111111;
	exp_table[11'b01111011110] = 16'b1111111111111111;
	exp_table[11'b01111011111] = 16'b1111111111111111;
	exp_table[11'b01111100000] = 16'b1111111111111111;
	exp_table[11'b01111100001] = 16'b1111111111111111;
	exp_table[11'b01111100010] = 16'b1111111111111111;
	exp_table[11'b01111100011] = 16'b1111111111111111;
	exp_table[11'b01111100100] = 16'b1111111111111111;
	exp_table[11'b01111100101] = 16'b1111111111111111;
	exp_table[11'b01111100110] = 16'b1111111111111111;
	exp_table[11'b01111100111] = 16'b1111111111111111;
	exp_table[11'b01111101000] = 16'b1111111111111111;
	exp_table[11'b01111101001] = 16'b1111111111111111;
	exp_table[11'b01111101010] = 16'b1111111111111111;
	exp_table[11'b01111101011] = 16'b1111111111111111;
	exp_table[11'b01111101100] = 16'b1111111111111111;
	exp_table[11'b01111101101] = 16'b1111111111111111;
	exp_table[11'b01111101110] = 16'b1111111111111111;
	exp_table[11'b01111101111] = 16'b1111111111111111;
	exp_table[11'b01111110000] = 16'b1111111111111111;
	exp_table[11'b01111110001] = 16'b1111111111111111;
	exp_table[11'b01111110010] = 16'b1111111111111111;
	exp_table[11'b01111110011] = 16'b1111111111111111;
	exp_table[11'b01111110100] = 16'b1111111111111111;
	exp_table[11'b01111110101] = 16'b1111111111111111;
	exp_table[11'b01111110110] = 16'b1111111111111111;
	exp_table[11'b01111110111] = 16'b1111111111111111;
	exp_table[11'b01111111000] = 16'b1111111111111111;
	exp_table[11'b01111111001] = 16'b1111111111111111;
	exp_table[11'b01111111010] = 16'b1111111111111111;
	exp_table[11'b01111111011] = 16'b1111111111111111;
	exp_table[11'b01111111100] = 16'b1111111111111111;
	exp_table[11'b01111111101] = 16'b1111111111111111;
	exp_table[11'b01111111110] = 16'b1111111111111111;
	exp_table[11'b01111111111] = 16'b1111111111111111;
    
    end
    
    always@(*)
    begin
        addr = in;
        exp_inner = exp_table[addr[16:6]];
    end
    
    assign exp = exp_inner;
endmodule